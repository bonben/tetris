--			when x"0001" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"0002" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"0003" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"0004" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"0005" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"0006" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"0007" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"0008" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"0009" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"000A" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"000B" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"000C" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"000D" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"000E" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"000F" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"0010" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"0011" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"0012" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"0013" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"0014" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"0015" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"0016" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"0017" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"0018" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"0019" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"001A" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"001B" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"001C" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"001D" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"001E" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"001F" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"0020" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"0021" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"0022" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"0023" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"0024" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"0025" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"0026" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"0027" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"0028" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"0029" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"002A" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"002B" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"002C" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"002D" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"002E" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"002F" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"0030" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"0031" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"0032" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"0033" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"0034" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"0035" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"0036" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"0037" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"0038" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"0039" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"003A" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"003B" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"003C" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"003D" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"003E" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"003F" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"0040" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"0041" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"0042" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"0043" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"0044" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"0045" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"0046" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"0047" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"0048" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"0049" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"004A" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"004B" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"004C" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"004D" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"004E" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"004F" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"0050" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"0051" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"0052" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"0053" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"0054" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"0055" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"0056" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"0057" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"0058" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"0059" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"005A" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"005B" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"005C" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"005D" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"005E" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"005F" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"0060" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"0061" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"0062" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"0063" => MILLIEMES <= x"0"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"0064" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"0065" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"0066" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"0067" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"0068" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"0069" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"006A" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"006B" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"006C" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"006D" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"006E" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"006F" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"0070" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"0071" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"0072" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"0073" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"0074" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"0075" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"0076" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"0077" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"0078" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"0079" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"007A" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"007B" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"007C" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"007D" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"007E" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"007F" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"0080" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"0081" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"0082" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"0083" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"0084" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"0085" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"0086" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"0087" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"0088" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"0089" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"008A" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"008B" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"008C" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"008D" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"008E" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"008F" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"0090" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"0091" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"0092" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"0093" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"0094" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"0095" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"0096" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"0097" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"0098" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"0099" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"009A" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"009B" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"009C" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"009D" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"009E" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"009F" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"00A0" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"00A1" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"00A2" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"00A3" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"00A4" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"00A5" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"00A6" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"00A7" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"00A8" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"00A9" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"00AA" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"00AB" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"00AC" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"00AD" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"00AE" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"00AF" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"00B0" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"00B1" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"00B2" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"00B3" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"00B4" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"00B5" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"00B6" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"00B7" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"00B8" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"00B9" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"00BA" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"00BB" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"00BC" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"00BD" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"00BE" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"00BF" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"00C0" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"00C1" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"00C2" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"00C3" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"00C4" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"00C5" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"00C6" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"00C7" => MILLIEMES <= x"0"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"00C8" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"00C9" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"00CA" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"00CB" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"00CC" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"00CD" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"00CE" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"00CF" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"00D0" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"00D1" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"00D2" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"00D3" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"00D4" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"00D5" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"00D6" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"00D7" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"00D8" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"00D9" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"00DA" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"00DB" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"00DC" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"00DD" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"00DE" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"00DF" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"00E0" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"00E1" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"00E2" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"00E3" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"00E4" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"00E5" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"00E6" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"00E7" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"00E8" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"00E9" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"00EA" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"00EB" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"00EC" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"00ED" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"00EE" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"00EF" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"00F0" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"00F1" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"00F2" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"00F3" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"00F4" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"00F5" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"00F6" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"00F7" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"00F8" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"00F9" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"00FA" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"00FB" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"00FC" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"00FD" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"00FE" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"00FF" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"0100" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"0101" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"0102" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"0103" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"0104" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"0105" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"0106" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"0107" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"0108" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"0109" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"010A" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"010B" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"010C" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"010D" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"010E" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"010F" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"0110" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"0111" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"0112" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"0113" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"0114" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"0115" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"0116" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"0117" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"0118" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"0119" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"011A" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"011B" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"011C" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"011D" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"011E" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"011F" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"0120" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"0121" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"0122" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"0123" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"0124" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"0125" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"0126" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"0127" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"0128" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"0129" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"012A" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"012B" => MILLIEMES <= x"0"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"012C" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"012D" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"012E" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"012F" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"0130" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"0131" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"0132" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"0133" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"0134" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"0135" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"0136" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"0137" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"0138" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"0139" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"013A" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"013B" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"013C" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"013D" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"013E" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"013F" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"0140" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"0141" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"0142" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"0143" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"0144" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"0145" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"0146" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"0147" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"0148" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"0149" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"014A" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"014B" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"014C" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"014D" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"014E" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"014F" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"0150" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"0151" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"0152" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"0153" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"0154" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"0155" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"0156" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"0157" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"0158" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"0159" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"015A" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"015B" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"015C" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"015D" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"015E" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"015F" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"0160" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"0161" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"0162" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"0163" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"0164" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"0165" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"0166" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"0167" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"0168" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"0169" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"016A" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"016B" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"016C" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"016D" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"016E" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"016F" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"0170" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"0171" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"0172" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"0173" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"0174" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"0175" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"0176" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"0177" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"0178" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"0179" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"017A" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"017B" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"017C" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"017D" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"017E" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"017F" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"0180" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"0181" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"0182" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"0183" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"0184" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"0185" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"0186" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"0187" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"0188" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"0189" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"018A" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"018B" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"018C" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"018D" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"018E" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"018F" => MILLIEMES <= x"0"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"0190" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"0191" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"0192" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"0193" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"0194" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"0195" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"0196" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"0197" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"0198" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"0199" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"019A" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"019B" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"019C" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"019D" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"019E" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"019F" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"01A0" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"01A1" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"01A2" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"01A3" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"01A4" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"01A5" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"01A6" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"01A7" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"01A8" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"01A9" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"01AA" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"01AB" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"01AC" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"01AD" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"01AE" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"01AF" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"01B0" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"01B1" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"01B2" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"01B3" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"01B4" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"01B5" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"01B6" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"01B7" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"01B8" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"01B9" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"01BA" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"01BB" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"01BC" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"01BD" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"01BE" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"01BF" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"01C0" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"01C1" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"01C2" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"01C3" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"01C4" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"01C5" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"01C6" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"01C7" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"01C8" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"01C9" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"01CA" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"01CB" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"01CC" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"01CD" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"01CE" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"01CF" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"01D0" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"01D1" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"01D2" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"01D3" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"01D4" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"01D5" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"01D6" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"01D7" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"01D8" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"01D9" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"01DA" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"01DB" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"01DC" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"01DD" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"01DE" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"01DF" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"01E0" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"01E1" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"01E2" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"01E3" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"01E4" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"01E5" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"01E6" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"01E7" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"01E8" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"01E9" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"01EA" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"01EB" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"01EC" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"01ED" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"01EE" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"01EF" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"01F0" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"01F1" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"01F2" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"01F3" => MILLIEMES <= x"0"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"01F4" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"01F5" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"01F6" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"01F7" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"01F8" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"01F9" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"01FA" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"01FB" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"01FC" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"01FD" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"01FE" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"01FF" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"0200" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"0201" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"0202" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"0203" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"0204" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"0205" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"0206" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"0207" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"0208" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"0209" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"020A" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"020B" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"020C" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"020D" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"020E" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"020F" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"0210" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"0211" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"0212" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"0213" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"0214" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"0215" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"0216" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"0217" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"0218" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"0219" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"021A" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"021B" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"021C" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"021D" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"021E" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"021F" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"0220" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"0221" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"0222" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"0223" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"0224" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"0225" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"0226" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"0227" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"0228" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"0229" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"022A" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"022B" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"022C" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"022D" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"022E" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"022F" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"0230" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"0231" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"0232" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"0233" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"0234" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"0235" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"0236" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"0237" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"0238" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"0239" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"023A" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"023B" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"023C" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"023D" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"023E" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"023F" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"0240" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"0241" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"0242" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"0243" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"0244" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"0245" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"0246" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"0247" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"0248" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"0249" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"024A" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"024B" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"024C" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"024D" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"024E" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"024F" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"0250" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"0251" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"0252" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"0253" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"0254" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"0255" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"0256" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"0257" => MILLIEMES <= x"0"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"0258" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"0259" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"025A" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"025B" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"025C" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"025D" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"025E" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"025F" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"0260" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"0261" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"0262" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"0263" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"0264" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"0265" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"0266" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"0267" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"0268" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"0269" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"026A" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"026B" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"026C" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"026D" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"026E" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"026F" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"0270" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"0271" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"0272" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"0273" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"0274" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"0275" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"0276" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"0277" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"0278" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"0279" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"027A" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"027B" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"027C" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"027D" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"027E" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"027F" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"0280" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"0281" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"0282" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"0283" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"0284" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"0285" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"0286" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"0287" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"0288" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"0289" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"028A" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"028B" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"028C" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"028D" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"028E" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"028F" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"0290" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"0291" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"0292" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"0293" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"0294" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"0295" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"0296" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"0297" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"0298" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"0299" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"029A" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"029B" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"029C" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"029D" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"029E" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"029F" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"02A0" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"02A1" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"02A2" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"02A3" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"02A4" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"02A5" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"02A6" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"02A7" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"02A8" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"02A9" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"02AA" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"02AB" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"02AC" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"02AD" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"02AE" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"02AF" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"02B0" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"02B1" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"02B2" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"02B3" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"02B4" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"02B5" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"02B6" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"02B7" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"02B8" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"02B9" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"02BA" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"02BB" => MILLIEMES <= x"0"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"02BC" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"02BD" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"02BE" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"02BF" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"02C0" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"02C1" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"02C2" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"02C3" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"02C4" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"02C5" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"02C6" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"02C7" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"02C8" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"02C9" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"02CA" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"02CB" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"02CC" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"02CD" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"02CE" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"02CF" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"02D0" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"02D1" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"02D2" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"02D3" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"02D4" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"02D5" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"02D6" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"02D7" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"02D8" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"02D9" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"02DA" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"02DB" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"02DC" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"02DD" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"02DE" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"02DF" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"02E0" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"02E1" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"02E2" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"02E3" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"02E4" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"02E5" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"02E6" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"02E7" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"02E8" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"02E9" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"02EA" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"02EB" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"02EC" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"02ED" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"02EE" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"02EF" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"02F0" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"02F1" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"02F2" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"02F3" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"02F4" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"02F5" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"02F6" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"02F7" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"02F8" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"02F9" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"02FA" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"02FB" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"02FC" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"02FD" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"02FE" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"02FF" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"0300" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"0301" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"0302" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"0303" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"0304" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"0305" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"0306" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"0307" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"0308" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"0309" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"030A" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"030B" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"030C" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"030D" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"030E" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"030F" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"0310" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"0311" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"0312" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"0313" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"0314" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"0315" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"0316" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"0317" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"0318" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"0319" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"031A" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"031B" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"031C" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"031D" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"031E" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"031F" => MILLIEMES <= x"0"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"0320" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"0321" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"0322" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"0323" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"0324" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"0325" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"0326" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"0327" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"0328" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"0329" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"032A" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"032B" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"032C" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"032D" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"032E" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"032F" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"0330" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"0331" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"0332" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"0333" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"0334" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"0335" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"0336" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"0337" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"0338" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"0339" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"033A" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"033B" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"033C" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"033D" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"033E" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"033F" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"0340" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"0341" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"0342" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"0343" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"0344" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"0345" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"0346" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"0347" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"0348" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"0349" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"034A" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"034B" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"034C" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"034D" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"034E" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"034F" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"0350" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"0351" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"0352" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"0353" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"0354" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"0355" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"0356" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"0357" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"0358" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"0359" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"035A" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"035B" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"035C" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"035D" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"035E" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"035F" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"0360" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"0361" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"0362" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"0363" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"0364" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"0365" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"0366" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"0367" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"0368" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"0369" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"036A" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"036B" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"036C" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"036D" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"036E" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"036F" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"0370" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"0371" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"0372" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"0373" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"0374" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"0375" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"0376" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"0377" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"0378" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"0379" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"037A" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"037B" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"037C" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"037D" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"037E" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"037F" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"0380" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"0381" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"0382" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"0383" => MILLIEMES <= x"0"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"0384" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"0385" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"0386" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"0387" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"0388" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"0389" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"038A" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"038B" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"038C" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"038D" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"038E" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"038F" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"0390" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"0391" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"0392" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"0393" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"0394" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"0395" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"0396" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"0397" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"0398" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"0399" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"039A" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"039B" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"039C" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"039D" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"039E" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"039F" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"03A0" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"03A1" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"03A2" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"03A3" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"03A4" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"03A5" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"03A6" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"03A7" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"03A8" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"03A9" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"03AA" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"03AB" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"03AC" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"03AD" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"03AE" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"03AF" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"03B0" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"03B1" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"03B2" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"03B3" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"03B4" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"03B5" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"03B6" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"03B7" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"03B8" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"03B9" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"03BA" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"03BB" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"03BC" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"03BD" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"03BE" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"03BF" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"03C0" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"03C1" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"03C2" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"03C3" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"03C4" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"03C5" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"03C6" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"03C7" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"03C8" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"03C9" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"03CA" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"03CB" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"03CC" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"03CD" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"03CE" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"03CF" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"03D0" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"03D1" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"03D2" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"03D3" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"03D4" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"03D5" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"03D6" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"03D7" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"03D8" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"03D9" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"03DA" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"03DB" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"03DC" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"03DD" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"03DE" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"03DF" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"03E0" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"03E1" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"03E2" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"03E3" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"03E4" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"03E5" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"03E6" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"03E7" => MILLIEMES <= x"0"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"03E8" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"03E9" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"03EA" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"03EB" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"03EC" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"03ED" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"03EE" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"03EF" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"03F0" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"03F1" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"03F2" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"03F3" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"03F4" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"03F5" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"03F6" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"03F7" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"03F8" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"03F9" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"03FA" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"03FB" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"03FC" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"03FD" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"03FE" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"03FF" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"0400" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"0401" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"0402" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"0403" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"0404" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"0405" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"0406" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"0407" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"0408" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"0409" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"040A" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"040B" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"040C" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"040D" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"040E" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"040F" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"0410" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"0411" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"0412" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"0413" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"0414" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"0415" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"0416" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"0417" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"0418" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"0419" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"041A" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"041B" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"041C" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"041D" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"041E" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"041F" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"0420" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"0421" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"0422" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"0423" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"0424" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"0425" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"0426" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"0427" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"0428" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"0429" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"042A" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"042B" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"042C" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"042D" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"042E" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"042F" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"0430" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"0431" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"0432" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"0433" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"0434" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"0435" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"0436" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"0437" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"0438" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"0439" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"043A" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"043B" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"043C" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"043D" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"043E" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"043F" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"0440" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"0441" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"0442" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"0443" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"0444" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"0445" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"0446" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"0447" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"0448" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"0449" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"044A" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"044B" => MILLIEMES <= x"1"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"044C" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"044D" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"044E" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"044F" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"0450" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"0451" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"0452" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"0453" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"0454" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"0455" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"0456" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"0457" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"0458" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"0459" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"045A" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"045B" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"045C" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"045D" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"045E" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"045F" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"0460" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"0461" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"0462" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"0463" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"0464" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"0465" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"0466" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"0467" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"0468" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"0469" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"046A" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"046B" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"046C" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"046D" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"046E" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"046F" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"0470" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"0471" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"0472" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"0473" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"0474" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"0475" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"0476" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"0477" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"0478" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"0479" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"047A" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"047B" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"047C" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"047D" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"047E" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"047F" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"0480" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"0481" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"0482" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"0483" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"0484" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"0485" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"0486" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"0487" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"0488" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"0489" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"048A" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"048B" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"048C" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"048D" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"048E" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"048F" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"0490" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"0491" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"0492" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"0493" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"0494" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"0495" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"0496" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"0497" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"0498" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"0499" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"049A" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"049B" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"049C" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"049D" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"049E" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"049F" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"04A0" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"04A1" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"04A2" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"04A3" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"04A4" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"04A5" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"04A6" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"04A7" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"04A8" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"04A9" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"04AA" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"04AB" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"04AC" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"04AD" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"04AE" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"04AF" => MILLIEMES <= x"1"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"04B0" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"04B1" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"04B2" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"04B3" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"04B4" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"04B5" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"04B6" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"04B7" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"04B8" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"04B9" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"04BA" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"04BB" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"04BC" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"04BD" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"04BE" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"04BF" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"04C0" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"04C1" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"04C2" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"04C3" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"04C4" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"04C5" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"04C6" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"04C7" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"04C8" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"04C9" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"04CA" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"04CB" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"04CC" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"04CD" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"04CE" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"04CF" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"04D0" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"04D1" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"04D2" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"04D3" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"04D4" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"04D5" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"04D6" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"04D7" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"04D8" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"04D9" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"04DA" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"04DB" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"04DC" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"04DD" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"04DE" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"04DF" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"04E0" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"04E1" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"04E2" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"04E3" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"04E4" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"04E5" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"04E6" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"04E7" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"04E8" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"04E9" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"04EA" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"04EB" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"04EC" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"04ED" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"04EE" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"04EF" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"04F0" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"04F1" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"04F2" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"04F3" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"04F4" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"04F5" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"04F6" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"04F7" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"04F8" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"04F9" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"04FA" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"04FB" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"04FC" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"04FD" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"04FE" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"04FF" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"0500" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"0501" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"0502" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"0503" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"0504" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"0505" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"0506" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"0507" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"0508" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"0509" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"050A" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"050B" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"050C" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"050D" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"050E" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"050F" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"0510" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"0511" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"0512" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"0513" => MILLIEMES <= x"1"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"0514" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"0515" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"0516" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"0517" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"0518" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"0519" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"051A" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"051B" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"051C" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"051D" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"051E" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"051F" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"0520" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"0521" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"0522" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"0523" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"0524" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"0525" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"0526" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"0527" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"0528" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"0529" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"052A" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"052B" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"052C" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"052D" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"052E" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"052F" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"0530" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"0531" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"0532" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"0533" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"0534" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"0535" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"0536" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"0537" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"0538" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"0539" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"053A" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"053B" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"053C" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"053D" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"053E" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"053F" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"0540" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"0541" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"0542" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"0543" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"0544" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"0545" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"0546" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"0547" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"0548" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"0549" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"054A" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"054B" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"054C" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"054D" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"054E" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"054F" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"0550" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"0551" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"0552" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"0553" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"0554" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"0555" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"0556" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"0557" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"0558" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"0559" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"055A" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"055B" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"055C" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"055D" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"055E" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"055F" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"0560" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"0561" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"0562" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"0563" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"0564" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"0565" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"0566" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"0567" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"0568" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"0569" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"056A" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"056B" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"056C" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"056D" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"056E" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"056F" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"0570" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"0571" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"0572" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"0573" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"0574" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"0575" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"0576" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"0577" => MILLIEMES <= x"1"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"0578" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"0579" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"057A" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"057B" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"057C" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"057D" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"057E" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"057F" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"0580" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"0581" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"0582" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"0583" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"0584" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"0585" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"0586" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"0587" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"0588" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"0589" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"058A" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"058B" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"058C" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"058D" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"058E" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"058F" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"0590" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"0591" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"0592" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"0593" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"0594" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"0595" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"0596" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"0597" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"0598" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"0599" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"059A" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"059B" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"059C" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"059D" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"059E" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"059F" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"05A0" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"05A1" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"05A2" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"05A3" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"05A4" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"05A5" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"05A6" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"05A7" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"05A8" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"05A9" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"05AA" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"05AB" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"05AC" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"05AD" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"05AE" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"05AF" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"05B0" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"05B1" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"05B2" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"05B3" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"05B4" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"05B5" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"05B6" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"05B7" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"05B8" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"05B9" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"05BA" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"05BB" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"05BC" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"05BD" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"05BE" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"05BF" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"05C0" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"05C1" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"05C2" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"05C3" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"05C4" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"05C5" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"05C6" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"05C7" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"05C8" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"05C9" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"05CA" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"05CB" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"05CC" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"05CD" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"05CE" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"05CF" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"05D0" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"05D1" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"05D2" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"05D3" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"05D4" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"05D5" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"05D6" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"05D7" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"05D8" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"05D9" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"05DA" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"05DB" => MILLIEMES <= x"1"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"05DC" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"05DD" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"05DE" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"05DF" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"05E0" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"05E1" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"05E2" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"05E3" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"05E4" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"05E5" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"05E6" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"05E7" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"05E8" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"05E9" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"05EA" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"05EB" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"05EC" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"05ED" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"05EE" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"05EF" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"05F0" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"05F1" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"05F2" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"05F3" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"05F4" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"05F5" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"05F6" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"05F7" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"05F8" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"05F9" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"05FA" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"05FB" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"05FC" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"05FD" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"05FE" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"05FF" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"0600" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"0601" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"0602" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"0603" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"0604" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"0605" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"0606" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"0607" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"0608" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"0609" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"060A" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"060B" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"060C" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"060D" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"060E" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"060F" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"0610" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"0611" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"0612" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"0613" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"0614" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"0615" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"0616" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"0617" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"0618" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"0619" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"061A" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"061B" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"061C" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"061D" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"061E" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"061F" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"0620" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"0621" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"0622" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"0623" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"0624" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"0625" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"0626" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"0627" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"0628" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"0629" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"062A" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"062B" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"062C" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"062D" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"062E" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"062F" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"0630" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"0631" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"0632" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"0633" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"0634" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"0635" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"0636" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"0637" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"0638" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"0639" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"063A" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"063B" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"063C" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"063D" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"063E" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"063F" => MILLIEMES <= x"1"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"0640" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"0641" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"0642" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"0643" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"0644" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"0645" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"0646" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"0647" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"0648" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"0649" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"064A" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"064B" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"064C" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"064D" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"064E" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"064F" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"0650" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"0651" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"0652" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"0653" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"0654" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"0655" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"0656" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"0657" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"0658" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"0659" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"065A" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"065B" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"065C" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"065D" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"065E" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"065F" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"0660" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"0661" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"0662" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"0663" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"0664" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"0665" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"0666" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"0667" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"0668" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"0669" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"066A" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"066B" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"066C" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"066D" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"066E" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"066F" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"0670" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"0671" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"0672" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"0673" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"0674" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"0675" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"0676" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"0677" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"0678" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"0679" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"067A" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"067B" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"067C" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"067D" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"067E" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"067F" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"0680" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"0681" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"0682" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"0683" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"0684" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"0685" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"0686" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"0687" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"0688" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"0689" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"068A" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"068B" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"068C" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"068D" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"068E" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"068F" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"0690" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"0691" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"0692" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"0693" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"0694" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"0695" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"0696" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"0697" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"0698" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"0699" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"069A" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"069B" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"069C" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"069D" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"069E" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"069F" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"06A0" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"06A1" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"06A2" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"06A3" => MILLIEMES <= x"1"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"06A4" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"06A5" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"06A6" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"06A7" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"06A8" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"06A9" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"06AA" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"06AB" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"06AC" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"06AD" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"06AE" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"06AF" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"06B0" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"06B1" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"06B2" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"06B3" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"06B4" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"06B5" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"06B6" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"06B7" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"06B8" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"06B9" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"06BA" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"06BB" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"06BC" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"06BD" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"06BE" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"06BF" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"06C0" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"06C1" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"06C2" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"06C3" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"06C4" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"06C5" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"06C6" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"06C7" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"06C8" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"06C9" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"06CA" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"06CB" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"06CC" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"06CD" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"06CE" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"06CF" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"06D0" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"06D1" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"06D2" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"06D3" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"06D4" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"06D5" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"06D6" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"06D7" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"06D8" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"06D9" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"06DA" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"06DB" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"06DC" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"06DD" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"06DE" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"06DF" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"06E0" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"06E1" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"06E2" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"06E3" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"06E4" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"06E5" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"06E6" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"06E7" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"06E8" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"06E9" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"06EA" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"06EB" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"06EC" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"06ED" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"06EE" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"06EF" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"06F0" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"06F1" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"06F2" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"06F3" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"06F4" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"06F5" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"06F6" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"06F7" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"06F8" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"06F9" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"06FA" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"06FB" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"06FC" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"06FD" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"06FE" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"06FF" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"0700" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"0701" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"0702" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"0703" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"0704" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"0705" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"0706" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"0707" => MILLIEMES <= x"1"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"0708" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"0709" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"070A" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"070B" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"070C" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"070D" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"070E" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"070F" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"0710" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"0711" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"0712" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"0713" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"0714" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"0715" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"0716" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"0717" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"0718" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"0719" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"071A" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"071B" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"071C" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"071D" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"071E" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"071F" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"0720" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"0721" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"0722" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"0723" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"0724" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"0725" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"0726" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"0727" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"0728" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"0729" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"072A" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"072B" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"072C" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"072D" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"072E" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"072F" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"0730" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"0731" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"0732" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"0733" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"0734" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"0735" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"0736" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"0737" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"0738" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"0739" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"073A" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"073B" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"073C" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"073D" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"073E" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"073F" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"0740" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"0741" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"0742" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"0743" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"0744" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"0745" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"0746" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"0747" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"0748" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"0749" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"074A" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"074B" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"074C" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"074D" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"074E" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"074F" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"0750" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"0751" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"0752" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"0753" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"0754" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"0755" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"0756" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"0757" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"0758" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"0759" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"075A" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"075B" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"075C" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"075D" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"075E" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"075F" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"0760" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"0761" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"0762" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"0763" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"0764" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"0765" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"0766" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"0767" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"0768" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"0769" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"076A" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"076B" => MILLIEMES <= x"1"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"076C" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"076D" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"076E" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"076F" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"0770" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"0771" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"0772" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"0773" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"0774" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"0775" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"0776" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"0777" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"0778" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"0779" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"077A" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"077B" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"077C" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"077D" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"077E" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"077F" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"0780" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"0781" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"0782" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"0783" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"0784" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"0785" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"0786" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"0787" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"0788" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"0789" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"078A" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"078B" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"078C" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"078D" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"078E" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"078F" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"0790" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"0791" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"0792" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"0793" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"0794" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"0795" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"0796" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"0797" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"0798" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"0799" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"079A" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"079B" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"079C" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"079D" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"079E" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"079F" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"07A0" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"07A1" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"07A2" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"07A3" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"07A4" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"07A5" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"07A6" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"07A7" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"07A8" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"07A9" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"07AA" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"07AB" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"07AC" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"07AD" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"07AE" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"07AF" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"07B0" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"07B1" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"07B2" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"07B3" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"07B4" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"07B5" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"07B6" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"07B7" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"07B8" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"07B9" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"07BA" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"07BB" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"07BC" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"07BD" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"07BE" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"07BF" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"07C0" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"07C1" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"07C2" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"07C3" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"07C4" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"07C5" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"07C6" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"07C7" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"07C8" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"07C9" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"07CA" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"07CB" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"07CC" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"07CD" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"07CE" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"07CF" => MILLIEMES <= x"1"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"07D0" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"07D1" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"07D2" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"07D3" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"07D4" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"07D5" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"07D6" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"07D7" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"07D8" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"07D9" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"07DA" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"07DB" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"07DC" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"07DD" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"07DE" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"07DF" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"07E0" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"07E1" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"07E2" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"07E3" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"07E4" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"07E5" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"07E6" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"07E7" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"07E8" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"07E9" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"07EA" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"07EB" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"07EC" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"07ED" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"07EE" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"07EF" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"07F0" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"07F1" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"07F2" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"07F3" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"07F4" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"07F5" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"07F6" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"07F7" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"07F8" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"07F9" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"07FA" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"07FB" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"07FC" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"07FD" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"07FE" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"07FF" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"0800" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"0801" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"0802" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"0803" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"0804" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"0805" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"0806" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"0807" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"0808" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"0809" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"080A" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"080B" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"080C" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"080D" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"080E" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"080F" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"0810" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"0811" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"0812" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"0813" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"0814" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"0815" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"0816" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"0817" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"0818" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"0819" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"081A" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"081B" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"081C" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"081D" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"081E" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"081F" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"0820" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"0821" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"0822" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"0823" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"0824" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"0825" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"0826" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"0827" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"0828" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"0829" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"082A" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"082B" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"082C" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"082D" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"082E" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"082F" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"0830" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"0831" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"0832" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"0833" => MILLIEMES <= x"2"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"0834" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"0835" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"0836" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"0837" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"0838" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"0839" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"083A" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"083B" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"083C" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"083D" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"083E" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"083F" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"0840" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"0841" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"0842" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"0843" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"0844" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"0845" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"0846" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"0847" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"0848" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"0849" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"084A" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"084B" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"084C" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"084D" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"084E" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"084F" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"0850" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"0851" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"0852" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"0853" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"0854" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"0855" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"0856" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"0857" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"0858" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"0859" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"085A" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"085B" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"085C" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"085D" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"085E" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"085F" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"0860" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"0861" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"0862" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"0863" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"0864" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"0865" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"0866" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"0867" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"0868" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"0869" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"086A" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"086B" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"086C" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"086D" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"086E" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"086F" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"0870" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"0871" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"0872" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"0873" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"0874" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"0875" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"0876" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"0877" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"0878" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"0879" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"087A" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"087B" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"087C" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"087D" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"087E" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"087F" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"0880" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"0881" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"0882" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"0883" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"0884" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"0885" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"0886" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"0887" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"0888" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"0889" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"088A" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"088B" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"088C" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"088D" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"088E" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"088F" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"0890" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"0891" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"0892" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"0893" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"0894" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"0895" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"0896" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"0897" => MILLIEMES <= x"2"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"0898" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"0899" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"089A" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"089B" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"089C" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"089D" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"089E" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"089F" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"08A0" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"08A1" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"08A2" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"08A3" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"08A4" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"08A5" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"08A6" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"08A7" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"08A8" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"08A9" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"08AA" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"08AB" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"08AC" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"08AD" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"08AE" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"08AF" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"08B0" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"08B1" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"08B2" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"08B3" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"08B4" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"08B5" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"08B6" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"08B7" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"08B8" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"08B9" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"08BA" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"08BB" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"08BC" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"08BD" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"08BE" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"08BF" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"08C0" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"08C1" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"08C2" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"08C3" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"08C4" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"08C5" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"08C6" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"08C7" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"08C8" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"08C9" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"08CA" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"08CB" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"08CC" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"08CD" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"08CE" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"08CF" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"08D0" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"08D1" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"08D2" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"08D3" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"08D4" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"08D5" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"08D6" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"08D7" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"08D8" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"08D9" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"08DA" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"08DB" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"08DC" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"08DD" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"08DE" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"08DF" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"08E0" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"08E1" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"08E2" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"08E3" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"08E4" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"08E5" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"08E6" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"08E7" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"08E8" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"08E9" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"08EA" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"08EB" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"08EC" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"08ED" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"08EE" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"08EF" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"08F0" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"08F1" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"08F2" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"08F3" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"08F4" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"08F5" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"08F6" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"08F7" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"08F8" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"08F9" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"08FA" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"08FB" => MILLIEMES <= x"2"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"08FC" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"08FD" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"08FE" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"08FF" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"0900" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"0901" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"0902" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"0903" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"0904" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"0905" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"0906" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"0907" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"0908" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"0909" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"090A" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"090B" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"090C" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"090D" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"090E" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"090F" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"0910" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"0911" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"0912" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"0913" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"0914" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"0915" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"0916" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"0917" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"0918" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"0919" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"091A" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"091B" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"091C" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"091D" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"091E" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"091F" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"0920" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"0921" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"0922" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"0923" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"0924" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"0925" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"0926" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"0927" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"0928" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"0929" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"092A" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"092B" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"092C" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"092D" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"092E" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"092F" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"0930" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"0931" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"0932" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"0933" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"0934" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"0935" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"0936" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"0937" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"0938" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"0939" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"093A" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"093B" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"093C" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"093D" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"093E" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"093F" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"0940" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"0941" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"0942" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"0943" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"0944" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"0945" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"0946" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"0947" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"0948" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"0949" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"094A" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"094B" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"094C" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"094D" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"094E" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"094F" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"0950" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"0951" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"0952" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"0953" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"0954" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"0955" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"0956" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"0957" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"0958" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"0959" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"095A" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"095B" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"095C" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"095D" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"095E" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"095F" => MILLIEMES <= x"2"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"0960" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"0961" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"0962" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"0963" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"0964" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"0965" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"0966" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"0967" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"0968" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"0969" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"096A" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"096B" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"096C" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"096D" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"096E" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"096F" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"0970" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"0971" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"0972" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"0973" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"0974" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"0975" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"0976" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"0977" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"0978" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"0979" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"097A" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"097B" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"097C" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"097D" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"097E" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"097F" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"0980" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"0981" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"0982" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"0983" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"0984" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"0985" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"0986" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"0987" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"0988" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"0989" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"098A" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"098B" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"098C" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"098D" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"098E" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"098F" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"0990" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"0991" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"0992" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"0993" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"0994" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"0995" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"0996" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"0997" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"0998" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"0999" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"099A" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"099B" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"099C" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"099D" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"099E" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"099F" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"09A0" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"09A1" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"09A2" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"09A3" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"09A4" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"09A5" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"09A6" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"09A7" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"09A8" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"09A9" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"09AA" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"09AB" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"09AC" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"09AD" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"09AE" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"09AF" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"09B0" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"09B1" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"09B2" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"09B3" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"09B4" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"09B5" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"09B6" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"09B7" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"09B8" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"09B9" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"09BA" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"09BB" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"09BC" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"09BD" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"09BE" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"09BF" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"09C0" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"09C1" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"09C2" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"09C3" => MILLIEMES <= x"2"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"09C4" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"09C5" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"09C6" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"09C7" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"09C8" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"09C9" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"09CA" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"09CB" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"09CC" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"09CD" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"09CE" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"09CF" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"09D0" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"09D1" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"09D2" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"09D3" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"09D4" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"09D5" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"09D6" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"09D7" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"09D8" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"09D9" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"09DA" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"09DB" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"09DC" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"09DD" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"09DE" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"09DF" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"09E0" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"09E1" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"09E2" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"09E3" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"09E4" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"09E5" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"09E6" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"09E7" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"09E8" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"09E9" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"09EA" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"09EB" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"09EC" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"09ED" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"09EE" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"09EF" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"09F0" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"09F1" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"09F2" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"09F3" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"09F4" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"09F5" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"09F6" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"09F7" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"09F8" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"09F9" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"09FA" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"09FB" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"09FC" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"09FD" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"09FE" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"09FF" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"0A00" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"0A01" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"0A02" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"0A03" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"0A04" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"0A05" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"0A06" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"0A07" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"0A08" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"0A09" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"0A0A" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"0A0B" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"0A0C" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"0A0D" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"0A0E" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"0A0F" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"0A10" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"0A11" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"0A12" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"0A13" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"0A14" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"0A15" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"0A16" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"0A17" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"0A18" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"0A19" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"0A1A" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"0A1B" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"0A1C" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"0A1D" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"0A1E" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"0A1F" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"0A20" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"0A21" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"0A22" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"0A23" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"0A24" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"0A25" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"0A26" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"0A27" => MILLIEMES <= x"2"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"0A28" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"0A29" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"0A2A" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"0A2B" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"0A2C" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"0A2D" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"0A2E" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"0A2F" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"0A30" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"0A31" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"0A32" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"0A33" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"0A34" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"0A35" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"0A36" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"0A37" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"0A38" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"0A39" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"0A3A" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"0A3B" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"0A3C" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"0A3D" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"0A3E" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"0A3F" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"0A40" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"0A41" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"0A42" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"0A43" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"0A44" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"0A45" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"0A46" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"0A47" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"0A48" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"0A49" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"0A4A" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"0A4B" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"0A4C" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"0A4D" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"0A4E" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"0A4F" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"0A50" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"0A51" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"0A52" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"0A53" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"0A54" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"0A55" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"0A56" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"0A57" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"0A58" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"0A59" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"0A5A" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"0A5B" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"0A5C" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"0A5D" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"0A5E" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"0A5F" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"0A60" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"0A61" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"0A62" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"0A63" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"0A64" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"0A65" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"0A66" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"0A67" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"0A68" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"0A69" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"0A6A" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"0A6B" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"0A6C" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"0A6D" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"0A6E" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"0A6F" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"0A70" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"0A71" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"0A72" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"0A73" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"0A74" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"0A75" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"0A76" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"0A77" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"0A78" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"0A79" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"0A7A" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"0A7B" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"0A7C" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"0A7D" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"0A7E" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"0A7F" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"0A80" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"0A81" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"0A82" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"0A83" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"0A84" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"0A85" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"0A86" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"0A87" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"0A88" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"0A89" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"0A8A" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"0A8B" => MILLIEMES <= x"2"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"0A8C" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"0A8D" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"0A8E" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"0A8F" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"0A90" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"0A91" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"0A92" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"0A93" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"0A94" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"0A95" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"0A96" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"0A97" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"0A98" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"0A99" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"0A9A" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"0A9B" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"0A9C" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"0A9D" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"0A9E" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"0A9F" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"0AA0" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"0AA1" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"0AA2" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"0AA3" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"0AA4" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"0AA5" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"0AA6" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"0AA7" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"0AA8" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"0AA9" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"0AAA" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"0AAB" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"0AAC" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"0AAD" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"0AAE" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"0AAF" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"0AB0" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"0AB1" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"0AB2" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"0AB3" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"0AB4" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"0AB5" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"0AB6" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"0AB7" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"0AB8" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"0AB9" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"0ABA" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"0ABB" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"0ABC" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"0ABD" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"0ABE" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"0ABF" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"0AC0" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"0AC1" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"0AC2" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"0AC3" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"0AC4" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"0AC5" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"0AC6" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"0AC7" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"0AC8" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"0AC9" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"0ACA" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"0ACB" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"0ACC" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"0ACD" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"0ACE" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"0ACF" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"0AD0" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"0AD1" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"0AD2" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"0AD3" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"0AD4" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"0AD5" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"0AD6" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"0AD7" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"0AD8" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"0AD9" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"0ADA" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"0ADB" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"0ADC" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"0ADD" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"0ADE" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"0ADF" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"0AE0" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"0AE1" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"0AE2" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"0AE3" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"0AE4" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"0AE5" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"0AE6" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"0AE7" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"0AE8" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"0AE9" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"0AEA" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"0AEB" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"0AEC" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"0AED" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"0AEE" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"0AEF" => MILLIEMES <= x"2"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"0AF0" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"0AF1" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"0AF2" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"0AF3" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"0AF4" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"0AF5" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"0AF6" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"0AF7" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"0AF8" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"0AF9" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"0AFA" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"0AFB" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"0AFC" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"0AFD" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"0AFE" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"0AFF" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"0B00" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"0B01" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"0B02" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"0B03" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"0B04" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"0B05" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"0B06" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"0B07" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"0B08" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"0B09" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"0B0A" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"0B0B" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"0B0C" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"0B0D" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"0B0E" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"0B0F" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"0B10" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"0B11" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"0B12" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"0B13" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"0B14" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"0B15" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"0B16" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"0B17" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"0B18" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"0B19" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"0B1A" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"0B1B" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"0B1C" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"0B1D" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"0B1E" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"0B1F" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"0B20" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"0B21" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"0B22" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"0B23" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"0B24" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"0B25" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"0B26" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"0B27" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"0B28" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"0B29" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"0B2A" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"0B2B" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"0B2C" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"0B2D" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"0B2E" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"0B2F" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"0B30" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"0B31" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"0B32" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"0B33" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"0B34" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"0B35" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"0B36" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"0B37" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"0B38" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"0B39" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"0B3A" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"0B3B" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"0B3C" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"0B3D" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"0B3E" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"0B3F" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"0B40" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"0B41" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"0B42" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"0B43" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"0B44" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"0B45" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"0B46" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"0B47" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"0B48" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"0B49" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"0B4A" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"0B4B" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"0B4C" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"0B4D" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"0B4E" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"0B4F" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"0B50" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"0B51" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"0B52" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"0B53" => MILLIEMES <= x"2"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"0B54" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"0B55" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"0B56" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"0B57" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"0B58" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"0B59" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"0B5A" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"0B5B" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"0B5C" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"0B5D" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"0B5E" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"0B5F" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"0B60" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"0B61" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"0B62" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"0B63" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"0B64" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"0B65" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"0B66" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"0B67" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"0B68" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"0B69" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"0B6A" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"0B6B" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"0B6C" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"0B6D" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"0B6E" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"0B6F" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"0B70" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"0B71" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"0B72" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"0B73" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"0B74" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"0B75" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"0B76" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"0B77" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"0B78" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"0B79" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"0B7A" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"0B7B" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"0B7C" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"0B7D" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"0B7E" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"0B7F" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"0B80" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"0B81" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"0B82" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"0B83" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"0B84" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"0B85" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"0B86" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"0B87" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"0B88" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"0B89" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"0B8A" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"0B8B" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"0B8C" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"0B8D" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"0B8E" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"0B8F" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"0B90" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"0B91" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"0B92" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"0B93" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"0B94" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"0B95" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"0B96" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"0B97" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"0B98" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"0B99" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"0B9A" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"0B9B" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"0B9C" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"0B9D" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"0B9E" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"0B9F" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"0BA0" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"0BA1" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"0BA2" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"0BA3" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"0BA4" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"0BA5" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"0BA6" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"0BA7" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"0BA8" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"0BA9" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"0BAA" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"0BAB" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"0BAC" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"0BAD" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"0BAE" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"0BAF" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"0BB0" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"0BB1" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"0BB2" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"0BB3" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"0BB4" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"0BB5" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"0BB6" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"0BB7" => MILLIEMES <= x"2"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"0BB8" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"0BB9" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"0BBA" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"0BBB" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"0BBC" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"0BBD" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"0BBE" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"0BBF" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"0BC0" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"0BC1" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"0BC2" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"0BC3" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"0BC4" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"0BC5" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"0BC6" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"0BC7" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"0BC8" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"0BC9" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"0BCA" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"0BCB" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"0BCC" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"0BCD" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"0BCE" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"0BCF" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"0BD0" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"0BD1" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"0BD2" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"0BD3" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"0BD4" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"0BD5" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"0BD6" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"0BD7" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"0BD8" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"0BD9" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"0BDA" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"0BDB" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"0BDC" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"0BDD" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"0BDE" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"0BDF" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"0BE0" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"0BE1" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"0BE2" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"0BE3" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"0BE4" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"0BE5" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"0BE6" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"0BE7" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"0BE8" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"0BE9" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"0BEA" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"0BEB" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"0BEC" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"0BED" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"0BEE" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"0BEF" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"0BF0" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"0BF1" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"0BF2" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"0BF3" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"0BF4" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"0BF5" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"0BF6" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"0BF7" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"0BF8" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"0BF9" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"0BFA" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"0BFB" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"0BFC" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"0BFD" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"0BFE" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"0BFF" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"0C00" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"0C01" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"0C02" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"0C03" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"0C04" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"0C05" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"0C06" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"0C07" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"0C08" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"0C09" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"0C0A" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"0C0B" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"0C0C" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"0C0D" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"0C0E" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"0C0F" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"0C10" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"0C11" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"0C12" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"0C13" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"0C14" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"0C15" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"0C16" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"0C17" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"0C18" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"0C19" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"0C1A" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"0C1B" => MILLIEMES <= x"3"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"0C1C" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"0C1D" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"0C1E" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"0C1F" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"0C20" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"0C21" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"0C22" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"0C23" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"0C24" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"0C25" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"0C26" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"0C27" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"0C28" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"0C29" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"0C2A" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"0C2B" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"0C2C" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"0C2D" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"0C2E" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"0C2F" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"0C30" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"0C31" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"0C32" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"0C33" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"0C34" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"0C35" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"0C36" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"0C37" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"0C38" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"0C39" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"0C3A" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"0C3B" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"0C3C" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"0C3D" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"0C3E" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"0C3F" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"0C40" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"0C41" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"0C42" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"0C43" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"0C44" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"0C45" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"0C46" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"0C47" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"0C48" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"0C49" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"0C4A" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"0C4B" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"0C4C" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"0C4D" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"0C4E" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"0C4F" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"0C50" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"0C51" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"0C52" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"0C53" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"0C54" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"0C55" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"0C56" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"0C57" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"0C58" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"0C59" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"0C5A" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"0C5B" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"0C5C" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"0C5D" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"0C5E" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"0C5F" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"0C60" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"0C61" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"0C62" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"0C63" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"0C64" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"0C65" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"0C66" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"0C67" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"0C68" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"0C69" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"0C6A" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"0C6B" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"0C6C" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"0C6D" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"0C6E" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"0C6F" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"0C70" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"0C71" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"0C72" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"0C73" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"0C74" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"0C75" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"0C76" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"0C77" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"0C78" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"0C79" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"0C7A" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"0C7B" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"0C7C" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"0C7D" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"0C7E" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"0C7F" => MILLIEMES <= x"3"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"0C80" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"0C81" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"0C82" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"0C83" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"0C84" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"0C85" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"0C86" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"0C87" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"0C88" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"0C89" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"0C8A" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"0C8B" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"0C8C" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"0C8D" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"0C8E" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"0C8F" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"0C90" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"0C91" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"0C92" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"0C93" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"0C94" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"0C95" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"0C96" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"0C97" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"0C98" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"0C99" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"0C9A" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"0C9B" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"0C9C" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"0C9D" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"0C9E" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"0C9F" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"0CA0" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"0CA1" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"0CA2" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"0CA3" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"0CA4" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"0CA5" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"0CA6" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"0CA7" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"0CA8" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"0CA9" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"0CAA" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"0CAB" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"0CAC" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"0CAD" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"0CAE" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"0CAF" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"0CB0" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"0CB1" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"0CB2" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"0CB3" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"0CB4" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"0CB5" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"0CB6" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"0CB7" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"0CB8" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"0CB9" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"0CBA" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"0CBB" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"0CBC" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"0CBD" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"0CBE" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"0CBF" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"0CC0" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"0CC1" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"0CC2" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"0CC3" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"0CC4" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"0CC5" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"0CC6" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"0CC7" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"0CC8" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"0CC9" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"0CCA" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"0CCB" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"0CCC" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"0CCD" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"0CCE" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"0CCF" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"0CD0" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"0CD1" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"0CD2" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"0CD3" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"0CD4" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"0CD5" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"0CD6" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"0CD7" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"0CD8" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"0CD9" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"0CDA" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"0CDB" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"0CDC" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"0CDD" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"0CDE" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"0CDF" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"0CE0" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"0CE1" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"0CE2" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"0CE3" => MILLIEMES <= x"3"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"0CE4" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"0CE5" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"0CE6" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"0CE7" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"0CE8" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"0CE9" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"0CEA" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"0CEB" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"0CEC" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"0CED" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"0CEE" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"0CEF" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"0CF0" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"0CF1" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"0CF2" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"0CF3" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"0CF4" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"0CF5" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"0CF6" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"0CF7" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"0CF8" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"0CF9" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"0CFA" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"0CFB" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"0CFC" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"0CFD" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"0CFE" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"0CFF" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"0D00" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"0D01" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"0D02" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"0D03" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"0D04" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"0D05" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"0D06" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"0D07" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"0D08" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"0D09" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"0D0A" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"0D0B" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"0D0C" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"0D0D" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"0D0E" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"0D0F" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"0D10" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"0D11" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"0D12" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"0D13" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"0D14" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"0D15" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"0D16" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"0D17" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"0D18" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"0D19" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"0D1A" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"0D1B" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"0D1C" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"0D1D" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"0D1E" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"0D1F" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"0D20" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"0D21" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"0D22" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"0D23" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"0D24" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"0D25" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"0D26" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"0D27" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"0D28" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"0D29" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"0D2A" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"0D2B" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"0D2C" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"0D2D" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"0D2E" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"0D2F" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"0D30" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"0D31" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"0D32" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"0D33" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"0D34" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"0D35" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"0D36" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"0D37" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"0D38" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"0D39" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"0D3A" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"0D3B" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"0D3C" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"0D3D" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"0D3E" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"0D3F" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"0D40" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"0D41" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"0D42" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"0D43" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"0D44" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"0D45" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"0D46" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"0D47" => MILLIEMES <= x"3"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"0D48" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"0D49" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"0D4A" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"0D4B" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"0D4C" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"0D4D" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"0D4E" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"0D4F" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"0D50" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"0D51" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"0D52" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"0D53" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"0D54" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"0D55" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"0D56" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"0D57" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"0D58" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"0D59" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"0D5A" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"0D5B" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"0D5C" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"0D5D" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"0D5E" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"0D5F" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"0D60" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"0D61" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"0D62" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"0D63" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"0D64" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"0D65" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"0D66" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"0D67" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"0D68" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"0D69" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"0D6A" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"0D6B" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"0D6C" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"0D6D" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"0D6E" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"0D6F" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"0D70" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"0D71" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"0D72" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"0D73" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"0D74" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"0D75" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"0D76" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"0D77" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"0D78" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"0D79" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"0D7A" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"0D7B" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"0D7C" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"0D7D" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"0D7E" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"0D7F" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"0D80" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"0D81" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"0D82" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"0D83" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"0D84" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"0D85" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"0D86" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"0D87" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"0D88" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"0D89" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"0D8A" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"0D8B" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"0D8C" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"0D8D" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"0D8E" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"0D8F" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"0D90" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"0D91" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"0D92" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"0D93" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"0D94" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"0D95" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"0D96" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"0D97" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"0D98" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"0D99" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"0D9A" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"0D9B" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"0D9C" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"0D9D" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"0D9E" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"0D9F" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"0DA0" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"0DA1" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"0DA2" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"0DA3" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"0DA4" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"0DA5" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"0DA6" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"0DA7" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"0DA8" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"0DA9" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"0DAA" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"0DAB" => MILLIEMES <= x"3"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"0DAC" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"0DAD" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"0DAE" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"0DAF" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"0DB0" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"0DB1" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"0DB2" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"0DB3" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"0DB4" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"0DB5" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"0DB6" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"0DB7" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"0DB8" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"0DB9" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"0DBA" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"0DBB" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"0DBC" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"0DBD" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"0DBE" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"0DBF" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"0DC0" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"0DC1" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"0DC2" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"0DC3" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"0DC4" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"0DC5" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"0DC6" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"0DC7" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"0DC8" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"0DC9" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"0DCA" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"0DCB" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"0DCC" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"0DCD" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"0DCE" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"0DCF" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"0DD0" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"0DD1" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"0DD2" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"0DD3" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"0DD4" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"0DD5" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"0DD6" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"0DD7" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"0DD8" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"0DD9" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"0DDA" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"0DDB" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"0DDC" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"0DDD" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"0DDE" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"0DDF" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"0DE0" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"0DE1" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"0DE2" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"0DE3" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"0DE4" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"0DE5" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"0DE6" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"0DE7" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"0DE8" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"0DE9" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"0DEA" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"0DEB" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"0DEC" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"0DED" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"0DEE" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"0DEF" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"0DF0" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"0DF1" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"0DF2" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"0DF3" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"0DF4" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"0DF5" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"0DF6" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"0DF7" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"0DF8" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"0DF9" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"0DFA" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"0DFB" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"0DFC" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"0DFD" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"0DFE" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"0DFF" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"0E00" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"0E01" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"0E02" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"0E03" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"0E04" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"0E05" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"0E06" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"0E07" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"0E08" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"0E09" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"0E0A" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"0E0B" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"0E0C" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"0E0D" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"0E0E" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"0E0F" => MILLIEMES <= x"3"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"0E10" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"0E11" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"0E12" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"0E13" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"0E14" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"0E15" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"0E16" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"0E17" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"0E18" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"0E19" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"0E1A" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"0E1B" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"0E1C" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"0E1D" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"0E1E" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"0E1F" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"0E20" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"0E21" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"0E22" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"0E23" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"0E24" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"0E25" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"0E26" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"0E27" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"0E28" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"0E29" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"0E2A" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"0E2B" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"0E2C" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"0E2D" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"0E2E" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"0E2F" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"0E30" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"0E31" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"0E32" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"0E33" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"0E34" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"0E35" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"0E36" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"0E37" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"0E38" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"0E39" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"0E3A" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"0E3B" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"0E3C" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"0E3D" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"0E3E" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"0E3F" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"0E40" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"0E41" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"0E42" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"0E43" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"0E44" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"0E45" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"0E46" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"0E47" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"0E48" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"0E49" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"0E4A" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"0E4B" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"0E4C" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"0E4D" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"0E4E" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"0E4F" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"0E50" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"0E51" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"0E52" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"0E53" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"0E54" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"0E55" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"0E56" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"0E57" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"0E58" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"0E59" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"0E5A" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"0E5B" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"0E5C" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"0E5D" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"0E5E" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"0E5F" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"0E60" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"0E61" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"0E62" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"0E63" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"0E64" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"0E65" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"0E66" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"0E67" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"0E68" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"0E69" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"0E6A" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"0E6B" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"0E6C" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"0E6D" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"0E6E" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"0E6F" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"0E70" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"0E71" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"0E72" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"0E73" => MILLIEMES <= x"3"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"0E74" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"0E75" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"0E76" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"0E77" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"0E78" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"0E79" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"0E7A" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"0E7B" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"0E7C" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"0E7D" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"0E7E" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"0E7F" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"0E80" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"0E81" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"0E82" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"0E83" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"0E84" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"0E85" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"0E86" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"0E87" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"0E88" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"0E89" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"0E8A" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"0E8B" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"0E8C" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"0E8D" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"0E8E" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"0E8F" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"0E90" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"0E91" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"0E92" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"0E93" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"0E94" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"0E95" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"0E96" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"0E97" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"0E98" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"0E99" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"0E9A" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"0E9B" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"0E9C" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"0E9D" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"0E9E" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"0E9F" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"0EA0" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"0EA1" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"0EA2" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"0EA3" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"0EA4" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"0EA5" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"0EA6" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"0EA7" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"0EA8" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"0EA9" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"0EAA" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"0EAB" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"0EAC" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"0EAD" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"0EAE" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"0EAF" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"0EB0" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"0EB1" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"0EB2" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"0EB3" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"0EB4" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"0EB5" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"0EB6" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"0EB7" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"0EB8" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"0EB9" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"0EBA" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"0EBB" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"0EBC" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"0EBD" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"0EBE" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"0EBF" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"0EC0" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"0EC1" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"0EC2" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"0EC3" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"0EC4" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"0EC5" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"0EC6" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"0EC7" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"0EC8" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"0EC9" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"0ECA" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"0ECB" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"0ECC" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"0ECD" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"0ECE" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"0ECF" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"0ED0" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"0ED1" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"0ED2" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"0ED3" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"0ED4" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"0ED5" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"0ED6" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"0ED7" => MILLIEMES <= x"3"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"0ED8" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"0ED9" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"0EDA" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"0EDB" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"0EDC" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"0EDD" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"0EDE" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"0EDF" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"0EE0" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"0EE1" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"0EE2" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"0EE3" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"0EE4" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"0EE5" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"0EE6" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"0EE7" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"0EE8" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"0EE9" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"0EEA" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"0EEB" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"0EEC" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"0EED" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"0EEE" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"0EEF" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"0EF0" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"0EF1" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"0EF2" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"0EF3" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"0EF4" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"0EF5" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"0EF6" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"0EF7" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"0EF8" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"0EF9" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"0EFA" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"0EFB" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"0EFC" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"0EFD" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"0EFE" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"0EFF" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"0F00" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"0F01" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"0F02" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"0F03" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"0F04" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"0F05" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"0F06" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"0F07" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"0F08" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"0F09" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"0F0A" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"0F0B" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"0F0C" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"0F0D" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"0F0E" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"0F0F" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"0F10" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"0F11" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"0F12" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"0F13" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"0F14" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"0F15" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"0F16" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"0F17" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"0F18" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"0F19" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"0F1A" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"0F1B" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"0F1C" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"0F1D" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"0F1E" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"0F1F" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"0F20" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"0F21" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"0F22" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"0F23" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"0F24" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"0F25" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"0F26" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"0F27" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"0F28" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"0F29" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"0F2A" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"0F2B" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"0F2C" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"0F2D" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"0F2E" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"0F2F" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"0F30" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"0F31" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"0F32" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"0F33" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"0F34" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"0F35" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"0F36" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"0F37" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"0F38" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"0F39" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"0F3A" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"0F3B" => MILLIEMES <= x"3"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"0F3C" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"0F3D" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"0F3E" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"0F3F" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"0F40" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"0F41" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"0F42" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"0F43" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"0F44" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"0F45" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"0F46" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"0F47" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"0F48" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"0F49" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"0F4A" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"0F4B" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"0F4C" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"0F4D" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"0F4E" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"0F4F" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"0F50" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"0F51" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"0F52" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"0F53" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"0F54" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"0F55" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"0F56" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"0F57" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"0F58" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"0F59" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"0F5A" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"0F5B" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"0F5C" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"0F5D" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"0F5E" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"0F5F" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"0F60" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"0F61" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"0F62" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"0F63" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"0F64" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"0F65" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"0F66" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"0F67" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"0F68" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"0F69" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"0F6A" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"0F6B" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"0F6C" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"0F6D" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"0F6E" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"0F6F" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"0F70" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"0F71" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"0F72" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"0F73" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"0F74" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"0F75" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"0F76" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"0F77" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"0F78" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"0F79" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"0F7A" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"0F7B" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"0F7C" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"0F7D" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"0F7E" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"0F7F" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"0F80" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"0F81" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"0F82" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"0F83" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"0F84" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"0F85" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"0F86" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"0F87" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"0F88" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"0F89" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"0F8A" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"0F8B" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"0F8C" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"0F8D" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"0F8E" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"0F8F" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"0F90" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"0F91" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"0F92" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"0F93" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"0F94" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"0F95" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"0F96" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"0F97" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"0F98" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"0F99" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"0F9A" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"0F9B" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"0F9C" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"0F9D" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"0F9E" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"0F9F" => MILLIEMES <= x"3"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"0FA0" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"0FA1" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"0FA2" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"0FA3" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"0FA4" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"0FA5" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"0FA6" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"0FA7" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"0FA8" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"0FA9" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"0FAA" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"0FAB" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"0FAC" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"0FAD" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"0FAE" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"0FAF" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"0FB0" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"0FB1" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"0FB2" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"0FB3" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"0FB4" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"0FB5" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"0FB6" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"0FB7" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"0FB8" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"0FB9" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"0FBA" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"0FBB" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"0FBC" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"0FBD" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"0FBE" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"0FBF" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"0FC0" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"0FC1" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"0FC2" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"0FC3" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"0FC4" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"0FC5" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"0FC6" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"0FC7" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"0FC8" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"0FC9" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"0FCA" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"0FCB" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"0FCC" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"0FCD" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"0FCE" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"0FCF" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"0FD0" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"0FD1" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"0FD2" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"0FD3" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"0FD4" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"0FD5" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"0FD6" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"0FD7" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"0FD8" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"0FD9" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"0FDA" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"0FDB" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"0FDC" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"0FDD" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"0FDE" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"0FDF" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"0FE0" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"0FE1" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"0FE2" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"0FE3" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"0FE4" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"0FE5" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"0FE6" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"0FE7" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"0FE8" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"0FE9" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"0FEA" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"0FEB" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"0FEC" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"0FED" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"0FEE" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"0FEF" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"0FF0" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"0FF1" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"0FF2" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"0FF3" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"0FF4" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"0FF5" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"0FF6" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"0FF7" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"0FF8" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"0FF9" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"0FFA" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"0FFB" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"0FFC" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"0FFD" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"0FFE" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"0FFF" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"1000" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"1001" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"1002" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"1003" => MILLIEMES <= x"4"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"1004" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"1005" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"1006" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"1007" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"1008" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"1009" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"100A" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"100B" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"100C" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"100D" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"100E" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"100F" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"1010" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"1011" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"1012" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"1013" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"1014" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"1015" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"1016" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"1017" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"1018" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"1019" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"101A" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"101B" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"101C" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"101D" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"101E" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"101F" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"1020" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"1021" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"1022" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"1023" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"1024" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"1025" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"1026" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"1027" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"1028" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"1029" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"102A" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"102B" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"102C" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"102D" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"102E" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"102F" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"1030" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"1031" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"1032" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"1033" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"1034" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"1035" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"1036" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"1037" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"1038" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"1039" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"103A" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"103B" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"103C" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"103D" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"103E" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"103F" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"1040" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"1041" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"1042" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"1043" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"1044" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"1045" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"1046" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"1047" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"1048" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"1049" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"104A" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"104B" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"104C" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"104D" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"104E" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"104F" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"1050" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"1051" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"1052" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"1053" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"1054" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"1055" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"1056" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"1057" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"1058" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"1059" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"105A" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"105B" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"105C" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"105D" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"105E" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"105F" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"1060" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"1061" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"1062" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"1063" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"1064" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"1065" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"1066" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"1067" => MILLIEMES <= x"4"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"1068" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"1069" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"106A" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"106B" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"106C" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"106D" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"106E" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"106F" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"1070" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"1071" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"1072" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"1073" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"1074" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"1075" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"1076" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"1077" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"1078" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"1079" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"107A" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"107B" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"107C" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"107D" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"107E" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"107F" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"1080" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"1081" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"1082" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"1083" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"1084" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"1085" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"1086" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"1087" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"1088" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"1089" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"108A" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"108B" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"108C" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"108D" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"108E" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"108F" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"1090" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"1091" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"1092" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"1093" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"1094" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"1095" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"1096" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"1097" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"1098" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"1099" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"109A" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"109B" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"109C" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"109D" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"109E" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"109F" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"10A0" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"10A1" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"10A2" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"10A3" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"10A4" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"10A5" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"10A6" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"10A7" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"10A8" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"10A9" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"10AA" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"10AB" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"10AC" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"10AD" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"10AE" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"10AF" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"10B0" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"10B1" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"10B2" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"10B3" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"10B4" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"10B5" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"10B6" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"10B7" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"10B8" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"10B9" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"10BA" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"10BB" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"10BC" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"10BD" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"10BE" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"10BF" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"10C0" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"10C1" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"10C2" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"10C3" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"10C4" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"10C5" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"10C6" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"10C7" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"10C8" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"10C9" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"10CA" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"10CB" => MILLIEMES <= x"4"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"10CC" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"10CD" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"10CE" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"10CF" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"10D0" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"10D1" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"10D2" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"10D3" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"10D4" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"10D5" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"10D6" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"10D7" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"10D8" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"10D9" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"10DA" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"10DB" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"10DC" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"10DD" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"10DE" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"10DF" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"10E0" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"10E1" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"10E2" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"10E3" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"10E4" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"10E5" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"10E6" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"10E7" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"10E8" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"10E9" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"10EA" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"10EB" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"10EC" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"10ED" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"10EE" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"10EF" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"10F0" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"10F1" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"10F2" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"10F3" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"10F4" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"10F5" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"10F6" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"10F7" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"10F8" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"10F9" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"10FA" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"10FB" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"10FC" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"10FD" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"10FE" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"10FF" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"1100" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"1101" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"1102" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"1103" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"1104" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"1105" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"1106" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"1107" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"1108" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"1109" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"110A" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"110B" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"110C" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"110D" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"110E" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"110F" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"1110" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"1111" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"1112" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"1113" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"1114" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"1115" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"1116" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"1117" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"1118" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"1119" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"111A" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"111B" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"111C" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"111D" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"111E" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"111F" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"1120" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"1121" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"1122" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"1123" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"1124" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"1125" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"1126" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"1127" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"1128" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"1129" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"112A" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"112B" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"112C" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"112D" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"112E" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"112F" => MILLIEMES <= x"4"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"1130" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"1131" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"1132" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"1133" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"1134" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"1135" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"1136" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"1137" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"1138" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"1139" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"113A" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"113B" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"113C" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"113D" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"113E" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"113F" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"1140" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"1141" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"1142" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"1143" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"1144" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"1145" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"1146" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"1147" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"1148" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"1149" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"114A" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"114B" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"114C" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"114D" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"114E" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"114F" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"1150" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"1151" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"1152" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"1153" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"1154" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"1155" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"1156" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"1157" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"1158" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"1159" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"115A" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"115B" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"115C" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"115D" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"115E" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"115F" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"1160" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"1161" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"1162" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"1163" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"1164" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"1165" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"1166" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"1167" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"1168" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"1169" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"116A" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"116B" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"116C" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"116D" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"116E" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"116F" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"1170" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"1171" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"1172" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"1173" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"1174" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"1175" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"1176" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"1177" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"1178" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"1179" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"117A" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"117B" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"117C" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"117D" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"117E" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"117F" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"1180" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"1181" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"1182" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"1183" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"1184" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"1185" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"1186" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"1187" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"1188" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"1189" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"118A" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"118B" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"118C" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"118D" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"118E" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"118F" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"1190" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"1191" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"1192" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"1193" => MILLIEMES <= x"4"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"1194" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"1195" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"1196" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"1197" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"1198" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"1199" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"119A" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"119B" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"119C" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"119D" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"119E" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"119F" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"11A0" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"11A1" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"11A2" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"11A3" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"11A4" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"11A5" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"11A6" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"11A7" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"11A8" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"11A9" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"11AA" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"11AB" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"11AC" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"11AD" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"11AE" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"11AF" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"11B0" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"11B1" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"11B2" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"11B3" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"11B4" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"11B5" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"11B6" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"11B7" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"11B8" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"11B9" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"11BA" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"11BB" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"11BC" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"11BD" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"11BE" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"11BF" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"11C0" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"11C1" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"11C2" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"11C3" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"11C4" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"11C5" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"11C6" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"11C7" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"11C8" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"11C9" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"11CA" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"11CB" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"11CC" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"11CD" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"11CE" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"11CF" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"11D0" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"11D1" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"11D2" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"11D3" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"11D4" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"11D5" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"11D6" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"11D7" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"11D8" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"11D9" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"11DA" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"11DB" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"11DC" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"11DD" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"11DE" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"11DF" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"11E0" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"11E1" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"11E2" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"11E3" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"11E4" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"11E5" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"11E6" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"11E7" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"11E8" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"11E9" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"11EA" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"11EB" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"11EC" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"11ED" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"11EE" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"11EF" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"11F0" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"11F1" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"11F2" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"11F3" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"11F4" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"11F5" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"11F6" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"11F7" => MILLIEMES <= x"4"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"11F8" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"11F9" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"11FA" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"11FB" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"11FC" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"11FD" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"11FE" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"11FF" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"1200" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"1201" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"1202" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"1203" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"1204" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"1205" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"1206" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"1207" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"1208" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"1209" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"120A" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"120B" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"120C" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"120D" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"120E" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"120F" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"1210" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"1211" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"1212" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"1213" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"1214" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"1215" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"1216" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"1217" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"1218" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"1219" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"121A" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"121B" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"121C" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"121D" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"121E" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"121F" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"1220" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"1221" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"1222" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"1223" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"1224" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"1225" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"1226" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"1227" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"1228" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"1229" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"122A" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"122B" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"122C" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"122D" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"122E" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"122F" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"1230" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"1231" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"1232" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"1233" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"1234" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"1235" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"1236" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"1237" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"1238" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"1239" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"123A" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"123B" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"123C" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"123D" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"123E" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"123F" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"1240" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"1241" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"1242" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"1243" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"1244" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"1245" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"1246" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"1247" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"1248" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"1249" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"124A" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"124B" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"124C" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"124D" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"124E" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"124F" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"1250" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"1251" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"1252" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"1253" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"1254" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"1255" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"1256" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"1257" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"1258" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"1259" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"125A" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"125B" => MILLIEMES <= x"4"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"125C" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"125D" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"125E" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"125F" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"1260" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"1261" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"1262" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"1263" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"1264" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"1265" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"1266" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"1267" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"1268" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"1269" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"126A" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"126B" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"126C" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"126D" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"126E" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"126F" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"1270" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"1271" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"1272" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"1273" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"1274" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"1275" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"1276" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"1277" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"1278" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"1279" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"127A" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"127B" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"127C" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"127D" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"127E" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"127F" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"1280" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"1281" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"1282" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"1283" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"1284" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"1285" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"1286" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"1287" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"1288" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"1289" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"128A" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"128B" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"128C" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"128D" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"128E" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"128F" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"1290" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"1291" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"1292" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"1293" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"1294" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"1295" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"1296" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"1297" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"1298" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"1299" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"129A" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"129B" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"129C" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"129D" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"129E" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"129F" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"12A0" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"12A1" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"12A2" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"12A3" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"12A4" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"12A5" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"12A6" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"12A7" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"12A8" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"12A9" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"12AA" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"12AB" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"12AC" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"12AD" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"12AE" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"12AF" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"12B0" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"12B1" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"12B2" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"12B3" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"12B4" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"12B5" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"12B6" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"12B7" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"12B8" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"12B9" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"12BA" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"12BB" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"12BC" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"12BD" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"12BE" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"12BF" => MILLIEMES <= x"4"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"12C0" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"12C1" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"12C2" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"12C3" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"12C4" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"12C5" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"12C6" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"12C7" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"12C8" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"12C9" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"12CA" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"12CB" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"12CC" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"12CD" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"12CE" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"12CF" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"12D0" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"12D1" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"12D2" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"12D3" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"12D4" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"12D5" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"12D6" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"12D7" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"12D8" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"12D9" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"12DA" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"12DB" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"12DC" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"12DD" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"12DE" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"12DF" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"12E0" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"12E1" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"12E2" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"12E3" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"12E4" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"12E5" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"12E6" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"12E7" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"12E8" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"12E9" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"12EA" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"12EB" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"12EC" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"12ED" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"12EE" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"12EF" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"12F0" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"12F1" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"12F2" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"12F3" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"12F4" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"12F5" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"12F6" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"12F7" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"12F8" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"12F9" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"12FA" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"12FB" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"12FC" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"12FD" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"12FE" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"12FF" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"1300" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"1301" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"1302" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"1303" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"1304" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"1305" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"1306" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"1307" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"1308" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"1309" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"130A" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"130B" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"130C" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"130D" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"130E" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"130F" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"1310" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"1311" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"1312" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"1313" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"1314" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"1315" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"1316" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"1317" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"1318" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"1319" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"131A" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"131B" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"131C" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"131D" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"131E" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"131F" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"1320" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"1321" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"1322" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"1323" => MILLIEMES <= x"4"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"1324" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"1325" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"1326" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"1327" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"1328" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"1329" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"132A" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"132B" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"132C" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"132D" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"132E" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"132F" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"1330" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"1331" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"1332" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"1333" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"1334" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"1335" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"1336" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"1337" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"1338" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"1339" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"133A" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"133B" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"133C" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"133D" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"133E" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"133F" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"1340" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"1341" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"1342" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"1343" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"1344" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"1345" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"1346" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"1347" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"1348" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"1349" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"134A" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"134B" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"134C" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"134D" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"134E" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"134F" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"1350" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"1351" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"1352" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"1353" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"1354" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"1355" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"1356" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"1357" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"1358" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"1359" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"135A" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"135B" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"135C" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"135D" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"135E" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"135F" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"1360" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"1361" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"1362" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"1363" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"1364" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"1365" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"1366" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"1367" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"1368" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"1369" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"136A" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"136B" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"136C" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"136D" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"136E" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"136F" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"1370" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"1371" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"1372" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"1373" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"1374" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"1375" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"1376" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"1377" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"1378" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"1379" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"137A" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"137B" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"137C" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"137D" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"137E" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"137F" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"1380" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"1381" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"1382" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"1383" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"1384" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"1385" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"1386" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"1387" => MILLIEMES <= x"4"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"1388" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"1389" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"138A" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"138B" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"138C" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"138D" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"138E" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"138F" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"1390" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"1391" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"1392" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"1393" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"1394" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"1395" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"1396" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"1397" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"1398" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"1399" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"139A" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"139B" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"139C" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"139D" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"139E" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"139F" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"13A0" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"13A1" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"13A2" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"13A3" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"13A4" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"13A5" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"13A6" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"13A7" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"13A8" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"13A9" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"13AA" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"13AB" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"13AC" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"13AD" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"13AE" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"13AF" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"13B0" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"13B1" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"13B2" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"13B3" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"13B4" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"13B5" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"13B6" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"13B7" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"13B8" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"13B9" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"13BA" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"13BB" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"13BC" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"13BD" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"13BE" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"13BF" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"13C0" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"13C1" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"13C2" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"13C3" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"13C4" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"13C5" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"13C6" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"13C7" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"13C8" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"13C9" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"13CA" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"13CB" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"13CC" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"13CD" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"13CE" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"13CF" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"13D0" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"13D1" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"13D2" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"13D3" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"13D4" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"13D5" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"13D6" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"13D7" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"13D8" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"13D9" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"13DA" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"13DB" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"13DC" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"13DD" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"13DE" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"13DF" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"13E0" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"13E1" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"13E2" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"13E3" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"13E4" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"13E5" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"13E6" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"13E7" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"13E8" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"13E9" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"13EA" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"13EB" => MILLIEMES <= x"5"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"13EC" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"13ED" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"13EE" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"13EF" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"13F0" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"13F1" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"13F2" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"13F3" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"13F4" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"13F5" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"13F6" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"13F7" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"13F8" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"13F9" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"13FA" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"13FB" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"13FC" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"13FD" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"13FE" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"13FF" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"1400" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"1401" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"1402" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"1403" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"1404" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"1405" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"1406" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"1407" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"1408" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"1409" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"140A" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"140B" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"140C" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"140D" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"140E" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"140F" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"1410" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"1411" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"1412" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"1413" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"1414" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"1415" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"1416" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"1417" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"1418" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"1419" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"141A" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"141B" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"141C" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"141D" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"141E" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"141F" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"1420" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"1421" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"1422" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"1423" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"1424" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"1425" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"1426" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"1427" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"1428" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"1429" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"142A" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"142B" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"142C" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"142D" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"142E" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"142F" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"1430" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"1431" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"1432" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"1433" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"1434" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"1435" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"1436" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"1437" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"1438" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"1439" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"143A" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"143B" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"143C" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"143D" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"143E" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"143F" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"1440" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"1441" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"1442" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"1443" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"1444" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"1445" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"1446" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"1447" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"1448" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"1449" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"144A" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"144B" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"144C" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"144D" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"144E" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"144F" => MILLIEMES <= x"5"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"1450" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"1451" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"1452" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"1453" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"1454" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"1455" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"1456" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"1457" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"1458" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"1459" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"145A" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"145B" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"145C" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"145D" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"145E" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"145F" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"1460" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"1461" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"1462" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"1463" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"1464" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"1465" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"1466" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"1467" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"1468" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"1469" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"146A" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"146B" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"146C" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"146D" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"146E" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"146F" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"1470" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"1471" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"1472" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"1473" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"1474" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"1475" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"1476" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"1477" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"1478" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"1479" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"147A" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"147B" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"147C" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"147D" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"147E" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"147F" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"1480" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"1481" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"1482" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"1483" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"1484" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"1485" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"1486" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"1487" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"1488" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"1489" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"148A" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"148B" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"148C" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"148D" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"148E" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"148F" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"1490" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"1491" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"1492" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"1493" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"1494" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"1495" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"1496" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"1497" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"1498" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"1499" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"149A" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"149B" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"149C" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"149D" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"149E" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"149F" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"14A0" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"14A1" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"14A2" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"14A3" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"14A4" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"14A5" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"14A6" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"14A7" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"14A8" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"14A9" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"14AA" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"14AB" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"14AC" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"14AD" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"14AE" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"14AF" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"14B0" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"14B1" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"14B2" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"14B3" => MILLIEMES <= x"5"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"14B4" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"14B5" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"14B6" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"14B7" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"14B8" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"14B9" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"14BA" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"14BB" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"14BC" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"14BD" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"14BE" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"14BF" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"14C0" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"14C1" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"14C2" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"14C3" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"14C4" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"14C5" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"14C6" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"14C7" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"14C8" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"14C9" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"14CA" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"14CB" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"14CC" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"14CD" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"14CE" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"14CF" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"14D0" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"14D1" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"14D2" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"14D3" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"14D4" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"14D5" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"14D6" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"14D7" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"14D8" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"14D9" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"14DA" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"14DB" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"14DC" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"14DD" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"14DE" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"14DF" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"14E0" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"14E1" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"14E2" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"14E3" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"14E4" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"14E5" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"14E6" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"14E7" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"14E8" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"14E9" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"14EA" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"14EB" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"14EC" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"14ED" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"14EE" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"14EF" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"14F0" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"14F1" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"14F2" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"14F3" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"14F4" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"14F5" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"14F6" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"14F7" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"14F8" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"14F9" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"14FA" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"14FB" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"14FC" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"14FD" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"14FE" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"14FF" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"1500" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"1501" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"1502" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"1503" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"1504" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"1505" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"1506" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"1507" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"1508" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"1509" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"150A" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"150B" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"150C" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"150D" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"150E" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"150F" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"1510" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"1511" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"1512" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"1513" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"1514" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"1515" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"1516" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"1517" => MILLIEMES <= x"5"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"1518" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"1519" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"151A" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"151B" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"151C" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"151D" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"151E" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"151F" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"1520" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"1521" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"1522" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"1523" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"1524" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"1525" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"1526" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"1527" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"1528" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"1529" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"152A" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"152B" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"152C" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"152D" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"152E" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"152F" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"1530" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"1531" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"1532" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"1533" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"1534" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"1535" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"1536" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"1537" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"1538" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"1539" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"153A" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"153B" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"153C" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"153D" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"153E" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"153F" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"1540" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"1541" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"1542" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"1543" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"1544" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"1545" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"1546" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"1547" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"1548" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"1549" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"154A" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"154B" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"154C" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"154D" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"154E" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"154F" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"1550" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"1551" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"1552" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"1553" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"1554" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"1555" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"1556" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"1557" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"1558" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"1559" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"155A" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"155B" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"155C" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"155D" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"155E" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"155F" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"1560" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"1561" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"1562" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"1563" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"1564" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"1565" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"1566" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"1567" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"1568" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"1569" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"156A" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"156B" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"156C" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"156D" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"156E" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"156F" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"1570" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"1571" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"1572" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"1573" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"1574" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"1575" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"1576" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"1577" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"1578" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"1579" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"157A" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"157B" => MILLIEMES <= x"5"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"157C" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"157D" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"157E" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"157F" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"1580" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"1581" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"1582" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"1583" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"1584" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"1585" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"1586" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"1587" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"1588" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"1589" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"158A" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"158B" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"158C" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"158D" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"158E" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"158F" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"1590" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"1591" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"1592" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"1593" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"1594" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"1595" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"1596" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"1597" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"1598" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"1599" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"159A" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"159B" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"159C" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"159D" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"159E" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"159F" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"15A0" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"15A1" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"15A2" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"15A3" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"15A4" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"15A5" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"15A6" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"15A7" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"15A8" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"15A9" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"15AA" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"15AB" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"15AC" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"15AD" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"15AE" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"15AF" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"15B0" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"15B1" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"15B2" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"15B3" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"15B4" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"15B5" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"15B6" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"15B7" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"15B8" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"15B9" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"15BA" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"15BB" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"15BC" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"15BD" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"15BE" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"15BF" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"15C0" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"15C1" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"15C2" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"15C3" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"15C4" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"15C5" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"15C6" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"15C7" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"15C8" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"15C9" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"15CA" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"15CB" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"15CC" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"15CD" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"15CE" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"15CF" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"15D0" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"15D1" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"15D2" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"15D3" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"15D4" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"15D5" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"15D6" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"15D7" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"15D8" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"15D9" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"15DA" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"15DB" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"15DC" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"15DD" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"15DE" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"15DF" => MILLIEMES <= x"5"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"15E0" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"15E1" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"15E2" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"15E3" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"15E4" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"15E5" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"15E6" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"15E7" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"15E8" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"15E9" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"15EA" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"15EB" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"15EC" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"15ED" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"15EE" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"15EF" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"15F0" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"15F1" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"15F2" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"15F3" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"15F4" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"15F5" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"15F6" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"15F7" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"15F8" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"15F9" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"15FA" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"15FB" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"15FC" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"15FD" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"15FE" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"15FF" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"1600" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"1601" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"1602" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"1603" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"1604" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"1605" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"1606" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"1607" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"1608" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"1609" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"160A" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"160B" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"160C" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"160D" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"160E" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"160F" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"1610" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"1611" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"1612" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"1613" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"1614" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"1615" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"1616" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"1617" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"1618" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"1619" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"161A" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"161B" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"161C" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"161D" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"161E" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"161F" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"1620" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"1621" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"1622" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"1623" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"1624" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"1625" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"1626" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"1627" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"1628" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"1629" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"162A" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"162B" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"162C" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"162D" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"162E" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"162F" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"1630" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"1631" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"1632" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"1633" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"1634" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"1635" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"1636" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"1637" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"1638" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"1639" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"163A" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"163B" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"163C" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"163D" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"163E" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"163F" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"1640" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"1641" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"1642" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"1643" => MILLIEMES <= x"5"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"1644" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"1645" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"1646" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"1647" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"1648" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"1649" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"164A" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"164B" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"164C" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"164D" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"164E" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"164F" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"1650" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"1651" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"1652" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"1653" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"1654" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"1655" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"1656" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"1657" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"1658" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"1659" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"165A" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"165B" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"165C" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"165D" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"165E" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"165F" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"1660" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"1661" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"1662" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"1663" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"1664" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"1665" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"1666" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"1667" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"1668" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"1669" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"166A" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"166B" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"166C" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"166D" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"166E" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"166F" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"1670" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"1671" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"1672" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"1673" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"1674" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"1675" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"1676" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"1677" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"1678" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"1679" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"167A" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"167B" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"167C" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"167D" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"167E" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"167F" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"1680" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"1681" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"1682" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"1683" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"1684" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"1685" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"1686" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"1687" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"1688" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"1689" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"168A" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"168B" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"168C" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"168D" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"168E" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"168F" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"1690" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"1691" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"1692" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"1693" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"1694" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"1695" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"1696" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"1697" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"1698" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"1699" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"169A" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"169B" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"169C" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"169D" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"169E" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"169F" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"16A0" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"16A1" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"16A2" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"16A3" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"16A4" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"16A5" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"16A6" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"16A7" => MILLIEMES <= x"5"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"16A8" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"16A9" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"16AA" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"16AB" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"16AC" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"16AD" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"16AE" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"16AF" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"16B0" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"16B1" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"16B2" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"16B3" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"16B4" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"16B5" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"16B6" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"16B7" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"16B8" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"16B9" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"16BA" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"16BB" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"16BC" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"16BD" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"16BE" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"16BF" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"16C0" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"16C1" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"16C2" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"16C3" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"16C4" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"16C5" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"16C6" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"16C7" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"16C8" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"16C9" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"16CA" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"16CB" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"16CC" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"16CD" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"16CE" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"16CF" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"16D0" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"16D1" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"16D2" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"16D3" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"16D4" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"16D5" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"16D6" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"16D7" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"16D8" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"16D9" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"16DA" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"16DB" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"16DC" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"16DD" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"16DE" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"16DF" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"16E0" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"16E1" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"16E2" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"16E3" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"16E4" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"16E5" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"16E6" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"16E7" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"16E8" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"16E9" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"16EA" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"16EB" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"16EC" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"16ED" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"16EE" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"16EF" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"16F0" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"16F1" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"16F2" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"16F3" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"16F4" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"16F5" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"16F6" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"16F7" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"16F8" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"16F9" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"16FA" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"16FB" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"16FC" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"16FD" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"16FE" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"16FF" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"1700" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"1701" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"1702" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"1703" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"1704" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"1705" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"1706" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"1707" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"1708" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"1709" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"170A" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"170B" => MILLIEMES <= x"5"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"170C" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"170D" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"170E" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"170F" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"1710" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"1711" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"1712" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"1713" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"1714" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"1715" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"1716" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"1717" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"1718" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"1719" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"171A" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"171B" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"171C" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"171D" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"171E" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"171F" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"1720" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"1721" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"1722" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"1723" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"1724" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"1725" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"1726" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"1727" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"1728" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"1729" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"172A" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"172B" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"172C" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"172D" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"172E" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"172F" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"1730" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"1731" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"1732" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"1733" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"1734" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"1735" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"1736" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"1737" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"1738" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"1739" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"173A" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"173B" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"173C" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"173D" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"173E" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"173F" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"1740" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"1741" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"1742" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"1743" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"1744" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"1745" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"1746" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"1747" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"1748" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"1749" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"174A" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"174B" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"174C" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"174D" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"174E" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"174F" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"1750" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"1751" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"1752" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"1753" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"1754" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"1755" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"1756" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"1757" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"1758" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"1759" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"175A" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"175B" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"175C" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"175D" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"175E" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"175F" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"1760" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"1761" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"1762" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"1763" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"1764" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"1765" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"1766" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"1767" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"1768" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"1769" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"176A" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"176B" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"176C" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"176D" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"176E" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"176F" => MILLIEMES <= x"5"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"1770" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"1771" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"1772" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"1773" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"1774" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"1775" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"1776" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"1777" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"1778" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"1779" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"177A" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"177B" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"177C" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"177D" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"177E" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"177F" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"1780" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"1781" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"1782" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"1783" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"1784" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"1785" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"1786" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"1787" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"1788" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"1789" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"178A" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"178B" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"178C" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"178D" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"178E" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"178F" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"1790" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"1791" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"1792" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"1793" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"1794" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"1795" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"1796" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"1797" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"1798" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"1799" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"179A" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"179B" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"179C" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"179D" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"179E" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"179F" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"17A0" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"17A1" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"17A2" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"17A3" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"17A4" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"17A5" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"17A6" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"17A7" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"17A8" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"17A9" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"17AA" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"17AB" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"17AC" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"17AD" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"17AE" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"17AF" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"17B0" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"17B1" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"17B2" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"17B3" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"17B4" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"17B5" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"17B6" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"17B7" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"17B8" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"17B9" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"17BA" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"17BB" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"17BC" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"17BD" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"17BE" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"17BF" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"17C0" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"17C1" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"17C2" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"17C3" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"17C4" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"17C5" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"17C6" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"17C7" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"17C8" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"17C9" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"17CA" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"17CB" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"17CC" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"17CD" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"17CE" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"17CF" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"17D0" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"17D1" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"17D2" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"17D3" => MILLIEMES <= x"6"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"17D4" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"17D5" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"17D6" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"17D7" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"17D8" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"17D9" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"17DA" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"17DB" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"17DC" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"17DD" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"17DE" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"17DF" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"17E0" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"17E1" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"17E2" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"17E3" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"17E4" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"17E5" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"17E6" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"17E7" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"17E8" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"17E9" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"17EA" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"17EB" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"17EC" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"17ED" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"17EE" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"17EF" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"17F0" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"17F1" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"17F2" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"17F3" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"17F4" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"17F5" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"17F6" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"17F7" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"17F8" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"17F9" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"17FA" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"17FB" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"17FC" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"17FD" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"17FE" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"17FF" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"1800" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"1801" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"1802" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"1803" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"1804" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"1805" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"1806" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"1807" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"1808" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"1809" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"180A" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"180B" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"180C" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"180D" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"180E" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"180F" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"1810" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"1811" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"1812" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"1813" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"1814" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"1815" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"1816" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"1817" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"1818" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"1819" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"181A" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"181B" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"181C" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"181D" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"181E" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"181F" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"1820" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"1821" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"1822" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"1823" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"1824" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"1825" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"1826" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"1827" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"1828" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"1829" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"182A" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"182B" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"182C" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"182D" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"182E" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"182F" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"1830" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"1831" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"1832" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"1833" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"1834" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"1835" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"1836" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"1837" => MILLIEMES <= x"6"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"1838" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"1839" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"183A" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"183B" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"183C" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"183D" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"183E" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"183F" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"1840" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"1841" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"1842" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"1843" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"1844" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"1845" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"1846" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"1847" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"1848" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"1849" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"184A" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"184B" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"184C" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"184D" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"184E" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"184F" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"1850" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"1851" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"1852" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"1853" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"1854" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"1855" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"1856" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"1857" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"1858" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"1859" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"185A" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"185B" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"185C" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"185D" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"185E" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"185F" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"1860" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"1861" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"1862" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"1863" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"1864" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"1865" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"1866" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"1867" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"1868" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"1869" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"186A" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"186B" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"186C" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"186D" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"186E" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"186F" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"1870" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"1871" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"1872" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"1873" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"1874" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"1875" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"1876" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"1877" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"1878" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"1879" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"187A" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"187B" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"187C" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"187D" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"187E" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"187F" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"1880" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"1881" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"1882" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"1883" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"1884" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"1885" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"1886" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"1887" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"1888" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"1889" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"188A" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"188B" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"188C" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"188D" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"188E" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"188F" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"1890" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"1891" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"1892" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"1893" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"1894" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"1895" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"1896" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"1897" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"1898" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"1899" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"189A" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"189B" => MILLIEMES <= x"6"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"189C" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"189D" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"189E" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"189F" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"18A0" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"18A1" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"18A2" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"18A3" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"18A4" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"18A5" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"18A6" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"18A7" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"18A8" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"18A9" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"18AA" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"18AB" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"18AC" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"18AD" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"18AE" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"18AF" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"18B0" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"18B1" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"18B2" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"18B3" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"18B4" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"18B5" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"18B6" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"18B7" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"18B8" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"18B9" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"18BA" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"18BB" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"18BC" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"18BD" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"18BE" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"18BF" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"18C0" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"18C1" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"18C2" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"18C3" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"18C4" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"18C5" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"18C6" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"18C7" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"18C8" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"18C9" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"18CA" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"18CB" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"18CC" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"18CD" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"18CE" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"18CF" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"18D0" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"18D1" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"18D2" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"18D3" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"18D4" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"18D5" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"18D6" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"18D7" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"18D8" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"18D9" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"18DA" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"18DB" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"18DC" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"18DD" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"18DE" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"18DF" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"18E0" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"18E1" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"18E2" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"18E3" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"18E4" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"18E5" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"18E6" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"18E7" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"18E8" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"18E9" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"18EA" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"18EB" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"18EC" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"18ED" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"18EE" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"18EF" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"18F0" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"18F1" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"18F2" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"18F3" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"18F4" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"18F5" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"18F6" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"18F7" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"18F8" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"18F9" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"18FA" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"18FB" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"18FC" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"18FD" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"18FE" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"18FF" => MILLIEMES <= x"6"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"1900" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"1901" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"1902" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"1903" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"1904" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"1905" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"1906" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"1907" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"1908" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"1909" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"190A" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"190B" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"190C" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"190D" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"190E" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"190F" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"1910" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"1911" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"1912" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"1913" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"1914" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"1915" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"1916" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"1917" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"1918" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"1919" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"191A" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"191B" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"191C" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"191D" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"191E" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"191F" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"1920" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"1921" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"1922" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"1923" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"1924" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"1925" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"1926" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"1927" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"1928" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"1929" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"192A" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"192B" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"192C" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"192D" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"192E" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"192F" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"1930" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"1931" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"1932" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"1933" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"1934" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"1935" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"1936" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"1937" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"1938" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"1939" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"193A" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"193B" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"193C" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"193D" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"193E" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"193F" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"1940" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"1941" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"1942" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"1943" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"1944" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"1945" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"1946" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"1947" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"1948" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"1949" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"194A" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"194B" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"194C" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"194D" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"194E" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"194F" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"1950" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"1951" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"1952" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"1953" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"1954" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"1955" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"1956" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"1957" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"1958" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"1959" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"195A" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"195B" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"195C" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"195D" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"195E" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"195F" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"1960" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"1961" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"1962" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"1963" => MILLIEMES <= x"6"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"1964" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"1965" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"1966" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"1967" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"1968" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"1969" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"196A" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"196B" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"196C" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"196D" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"196E" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"196F" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"1970" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"1971" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"1972" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"1973" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"1974" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"1975" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"1976" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"1977" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"1978" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"1979" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"197A" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"197B" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"197C" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"197D" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"197E" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"197F" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"1980" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"1981" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"1982" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"1983" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"1984" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"1985" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"1986" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"1987" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"1988" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"1989" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"198A" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"198B" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"198C" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"198D" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"198E" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"198F" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"1990" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"1991" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"1992" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"1993" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"1994" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"1995" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"1996" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"1997" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"1998" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"1999" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"199A" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"199B" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"199C" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"199D" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"199E" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"199F" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"19A0" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"19A1" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"19A2" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"19A3" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"19A4" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"19A5" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"19A6" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"19A7" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"19A8" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"19A9" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"19AA" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"19AB" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"19AC" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"19AD" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"19AE" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"19AF" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"19B0" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"19B1" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"19B2" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"19B3" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"19B4" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"19B5" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"19B6" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"19B7" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"19B8" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"19B9" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"19BA" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"19BB" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"19BC" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"19BD" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"19BE" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"19BF" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"19C0" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"19C1" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"19C2" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"19C3" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"19C4" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"19C5" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"19C6" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"19C7" => MILLIEMES <= x"6"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"19C8" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"19C9" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"19CA" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"19CB" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"19CC" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"19CD" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"19CE" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"19CF" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"19D0" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"19D1" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"19D2" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"19D3" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"19D4" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"19D5" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"19D6" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"19D7" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"19D8" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"19D9" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"19DA" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"19DB" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"19DC" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"19DD" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"19DE" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"19DF" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"19E0" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"19E1" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"19E2" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"19E3" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"19E4" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"19E5" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"19E6" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"19E7" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"19E8" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"19E9" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"19EA" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"19EB" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"19EC" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"19ED" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"19EE" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"19EF" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"19F0" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"19F1" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"19F2" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"19F3" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"19F4" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"19F5" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"19F6" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"19F7" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"19F8" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"19F9" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"19FA" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"19FB" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"19FC" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"19FD" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"19FE" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"19FF" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"1A00" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"1A01" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"1A02" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"1A03" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"1A04" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"1A05" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"1A06" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"1A07" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"1A08" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"1A09" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"1A0A" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"1A0B" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"1A0C" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"1A0D" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"1A0E" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"1A0F" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"1A10" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"1A11" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"1A12" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"1A13" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"1A14" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"1A15" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"1A16" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"1A17" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"1A18" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"1A19" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"1A1A" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"1A1B" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"1A1C" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"1A1D" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"1A1E" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"1A1F" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"1A20" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"1A21" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"1A22" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"1A23" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"1A24" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"1A25" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"1A26" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"1A27" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"1A28" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"1A29" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"1A2A" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"1A2B" => MILLIEMES <= x"6"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"1A2C" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"1A2D" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"1A2E" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"1A2F" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"1A30" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"1A31" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"1A32" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"1A33" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"1A34" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"1A35" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"1A36" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"1A37" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"1A38" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"1A39" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"1A3A" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"1A3B" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"1A3C" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"1A3D" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"1A3E" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"1A3F" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"1A40" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"1A41" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"1A42" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"1A43" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"1A44" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"1A45" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"1A46" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"1A47" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"1A48" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"1A49" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"1A4A" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"1A4B" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"1A4C" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"1A4D" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"1A4E" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"1A4F" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"1A50" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"1A51" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"1A52" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"1A53" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"1A54" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"1A55" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"1A56" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"1A57" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"1A58" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"1A59" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"1A5A" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"1A5B" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"1A5C" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"1A5D" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"1A5E" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"1A5F" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"1A60" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"1A61" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"1A62" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"1A63" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"1A64" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"1A65" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"1A66" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"1A67" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"1A68" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"1A69" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"1A6A" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"1A6B" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"1A6C" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"1A6D" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"1A6E" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"1A6F" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"1A70" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"1A71" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"1A72" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"1A73" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"1A74" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"1A75" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"1A76" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"1A77" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"1A78" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"1A79" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"1A7A" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"1A7B" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"1A7C" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"1A7D" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"1A7E" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"1A7F" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"1A80" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"1A81" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"1A82" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"1A83" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"1A84" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"1A85" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"1A86" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"1A87" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"1A88" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"1A89" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"1A8A" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"1A8B" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"1A8C" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"1A8D" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"1A8E" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"1A8F" => MILLIEMES <= x"6"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"1A90" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"1A91" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"1A92" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"1A93" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"1A94" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"1A95" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"1A96" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"1A97" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"1A98" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"1A99" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"1A9A" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"1A9B" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"1A9C" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"1A9D" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"1A9E" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"1A9F" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"1AA0" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"1AA1" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"1AA2" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"1AA3" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"1AA4" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"1AA5" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"1AA6" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"1AA7" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"1AA8" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"1AA9" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"1AAA" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"1AAB" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"1AAC" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"1AAD" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"1AAE" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"1AAF" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"1AB0" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"1AB1" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"1AB2" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"1AB3" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"1AB4" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"1AB5" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"1AB6" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"1AB7" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"1AB8" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"1AB9" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"1ABA" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"1ABB" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"1ABC" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"1ABD" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"1ABE" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"1ABF" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"1AC0" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"1AC1" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"1AC2" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"1AC3" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"1AC4" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"1AC5" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"1AC6" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"1AC7" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"1AC8" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"1AC9" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"1ACA" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"1ACB" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"1ACC" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"1ACD" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"1ACE" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"1ACF" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"1AD0" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"1AD1" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"1AD2" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"1AD3" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"1AD4" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"1AD5" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"1AD6" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"1AD7" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"1AD8" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"1AD9" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"1ADA" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"1ADB" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"1ADC" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"1ADD" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"1ADE" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"1ADF" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"1AE0" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"1AE1" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"1AE2" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"1AE3" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"1AE4" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"1AE5" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"1AE6" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"1AE7" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"1AE8" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"1AE9" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"1AEA" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"1AEB" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"1AEC" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"1AED" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"1AEE" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"1AEF" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"1AF0" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"1AF1" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"1AF2" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"1AF3" => MILLIEMES <= x"6"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"1AF4" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"1AF5" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"1AF6" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"1AF7" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"1AF8" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"1AF9" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"1AFA" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"1AFB" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"1AFC" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"1AFD" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"1AFE" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"1AFF" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"1B00" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"1B01" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"1B02" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"1B03" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"1B04" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"1B05" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"1B06" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"1B07" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"1B08" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"1B09" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"1B0A" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"1B0B" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"1B0C" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"1B0D" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"1B0E" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"1B0F" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"1B10" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"1B11" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"1B12" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"1B13" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"1B14" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"1B15" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"1B16" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"1B17" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"1B18" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"1B19" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"1B1A" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"1B1B" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"1B1C" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"1B1D" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"1B1E" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"1B1F" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"1B20" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"1B21" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"1B22" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"1B23" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"1B24" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"1B25" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"1B26" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"1B27" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"1B28" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"1B29" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"1B2A" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"1B2B" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"1B2C" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"1B2D" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"1B2E" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"1B2F" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"1B30" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"1B31" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"1B32" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"1B33" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"1B34" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"1B35" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"1B36" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"1B37" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"1B38" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"1B39" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"1B3A" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"1B3B" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"1B3C" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"1B3D" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"1B3E" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"1B3F" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"1B40" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"1B41" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"1B42" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"1B43" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"1B44" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"1B45" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"1B46" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"1B47" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"1B48" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"1B49" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"1B4A" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"1B4B" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"1B4C" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"1B4D" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"1B4E" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"1B4F" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"1B50" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"1B51" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"1B52" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"1B53" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"1B54" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"1B55" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"1B56" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"1B57" => MILLIEMES <= x"6"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"1B58" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"1B59" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"1B5A" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"1B5B" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"1B5C" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"1B5D" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"1B5E" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"1B5F" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"1B60" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"1B61" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"1B62" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"1B63" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"1B64" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"1B65" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"1B66" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"1B67" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"1B68" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"1B69" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"1B6A" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"1B6B" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"1B6C" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"1B6D" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"1B6E" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"1B6F" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"1B70" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"1B71" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"1B72" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"1B73" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"1B74" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"1B75" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"1B76" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"1B77" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"1B78" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"1B79" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"1B7A" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"1B7B" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"1B7C" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"1B7D" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"1B7E" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"1B7F" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"1B80" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"1B81" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"1B82" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"1B83" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"1B84" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"1B85" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"1B86" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"1B87" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"1B88" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"1B89" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"1B8A" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"1B8B" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"1B8C" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"1B8D" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"1B8E" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"1B8F" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"1B90" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"1B91" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"1B92" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"1B93" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"1B94" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"1B95" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"1B96" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"1B97" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"1B98" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"1B99" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"1B9A" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"1B9B" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"1B9C" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"1B9D" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"1B9E" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"1B9F" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"1BA0" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"1BA1" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"1BA2" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"1BA3" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"1BA4" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"1BA5" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"1BA6" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"1BA7" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"1BA8" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"1BA9" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"1BAA" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"1BAB" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"1BAC" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"1BAD" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"1BAE" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"1BAF" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"1BB0" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"1BB1" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"1BB2" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"1BB3" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"1BB4" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"1BB5" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"1BB6" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"1BB7" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"1BB8" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"1BB9" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"1BBA" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"1BBB" => MILLIEMES <= x"7"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"1BBC" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"1BBD" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"1BBE" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"1BBF" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"1BC0" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"1BC1" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"1BC2" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"1BC3" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"1BC4" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"1BC5" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"1BC6" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"1BC7" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"1BC8" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"1BC9" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"1BCA" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"1BCB" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"1BCC" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"1BCD" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"1BCE" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"1BCF" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"1BD0" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"1BD1" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"1BD2" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"1BD3" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"1BD4" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"1BD5" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"1BD6" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"1BD7" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"1BD8" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"1BD9" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"1BDA" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"1BDB" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"1BDC" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"1BDD" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"1BDE" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"1BDF" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"1BE0" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"1BE1" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"1BE2" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"1BE3" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"1BE4" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"1BE5" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"1BE6" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"1BE7" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"1BE8" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"1BE9" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"1BEA" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"1BEB" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"1BEC" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"1BED" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"1BEE" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"1BEF" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"1BF0" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"1BF1" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"1BF2" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"1BF3" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"1BF4" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"1BF5" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"1BF6" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"1BF7" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"1BF8" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"1BF9" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"1BFA" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"1BFB" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"1BFC" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"1BFD" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"1BFE" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"1BFF" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"1C00" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"1C01" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"1C02" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"1C03" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"1C04" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"1C05" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"1C06" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"1C07" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"1C08" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"1C09" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"1C0A" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"1C0B" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"1C0C" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"1C0D" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"1C0E" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"1C0F" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"1C10" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"1C11" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"1C12" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"1C13" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"1C14" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"1C15" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"1C16" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"1C17" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"1C18" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"1C19" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"1C1A" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"1C1B" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"1C1C" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"1C1D" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"1C1E" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"1C1F" => MILLIEMES <= x"7"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"1C20" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"1C21" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"1C22" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"1C23" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"1C24" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"1C25" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"1C26" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"1C27" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"1C28" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"1C29" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"1C2A" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"1C2B" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"1C2C" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"1C2D" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"1C2E" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"1C2F" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"1C30" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"1C31" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"1C32" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"1C33" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"1C34" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"1C35" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"1C36" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"1C37" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"1C38" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"1C39" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"1C3A" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"1C3B" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"1C3C" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"1C3D" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"1C3E" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"1C3F" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"1C40" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"1C41" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"1C42" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"1C43" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"1C44" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"1C45" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"1C46" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"1C47" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"1C48" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"1C49" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"1C4A" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"1C4B" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"1C4C" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"1C4D" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"1C4E" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"1C4F" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"1C50" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"1C51" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"1C52" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"1C53" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"1C54" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"1C55" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"1C56" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"1C57" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"1C58" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"1C59" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"1C5A" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"1C5B" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"1C5C" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"1C5D" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"1C5E" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"1C5F" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"1C60" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"1C61" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"1C62" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"1C63" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"1C64" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"1C65" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"1C66" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"1C67" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"1C68" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"1C69" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"1C6A" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"1C6B" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"1C6C" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"1C6D" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"1C6E" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"1C6F" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"1C70" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"1C71" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"1C72" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"1C73" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"1C74" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"1C75" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"1C76" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"1C77" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"1C78" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"1C79" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"1C7A" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"1C7B" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"1C7C" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"1C7D" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"1C7E" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"1C7F" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"1C80" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"1C81" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"1C82" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"1C83" => MILLIEMES <= x"7"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"1C84" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"1C85" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"1C86" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"1C87" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"1C88" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"1C89" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"1C8A" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"1C8B" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"1C8C" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"1C8D" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"1C8E" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"1C8F" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"1C90" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"1C91" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"1C92" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"1C93" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"1C94" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"1C95" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"1C96" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"1C97" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"1C98" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"1C99" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"1C9A" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"1C9B" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"1C9C" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"1C9D" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"1C9E" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"1C9F" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"1CA0" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"1CA1" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"1CA2" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"1CA3" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"1CA4" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"1CA5" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"1CA6" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"1CA7" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"1CA8" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"1CA9" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"1CAA" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"1CAB" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"1CAC" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"1CAD" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"1CAE" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"1CAF" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"1CB0" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"1CB1" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"1CB2" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"1CB3" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"1CB4" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"1CB5" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"1CB6" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"1CB7" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"1CB8" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"1CB9" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"1CBA" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"1CBB" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"1CBC" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"1CBD" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"1CBE" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"1CBF" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"1CC0" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"1CC1" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"1CC2" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"1CC3" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"1CC4" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"1CC5" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"1CC6" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"1CC7" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"1CC8" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"1CC9" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"1CCA" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"1CCB" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"1CCC" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"1CCD" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"1CCE" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"1CCF" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"1CD0" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"1CD1" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"1CD2" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"1CD3" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"1CD4" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"1CD5" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"1CD6" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"1CD7" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"1CD8" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"1CD9" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"1CDA" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"1CDB" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"1CDC" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"1CDD" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"1CDE" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"1CDF" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"1CE0" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"1CE1" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"1CE2" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"1CE3" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"1CE4" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"1CE5" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"1CE6" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"1CE7" => MILLIEMES <= x"7"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"1CE8" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"1CE9" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"1CEA" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"1CEB" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"1CEC" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"1CED" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"1CEE" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"1CEF" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"1CF0" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"1CF1" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"1CF2" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"1CF3" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"1CF4" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"1CF5" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"1CF6" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"1CF7" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"1CF8" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"1CF9" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"1CFA" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"1CFB" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"1CFC" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"1CFD" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"1CFE" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"1CFF" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"1D00" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"1D01" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"1D02" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"1D03" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"1D04" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"1D05" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"1D06" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"1D07" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"1D08" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"1D09" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"1D0A" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"1D0B" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"1D0C" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"1D0D" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"1D0E" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"1D0F" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"1D10" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"1D11" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"1D12" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"1D13" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"1D14" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"1D15" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"1D16" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"1D17" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"1D18" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"1D19" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"1D1A" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"1D1B" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"1D1C" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"1D1D" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"1D1E" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"1D1F" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"1D20" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"1D21" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"1D22" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"1D23" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"1D24" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"1D25" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"1D26" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"1D27" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"1D28" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"1D29" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"1D2A" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"1D2B" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"1D2C" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"1D2D" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"1D2E" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"1D2F" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"1D30" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"1D31" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"1D32" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"1D33" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"1D34" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"1D35" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"1D36" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"1D37" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"1D38" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"1D39" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"1D3A" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"1D3B" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"1D3C" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"1D3D" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"1D3E" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"1D3F" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"1D40" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"1D41" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"1D42" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"1D43" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"1D44" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"1D45" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"1D46" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"1D47" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"1D48" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"1D49" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"1D4A" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"1D4B" => MILLIEMES <= x"7"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"1D4C" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"1D4D" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"1D4E" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"1D4F" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"1D50" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"1D51" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"1D52" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"1D53" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"1D54" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"1D55" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"1D56" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"1D57" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"1D58" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"1D59" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"1D5A" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"1D5B" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"1D5C" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"1D5D" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"1D5E" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"1D5F" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"1D60" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"1D61" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"1D62" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"1D63" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"1D64" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"1D65" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"1D66" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"1D67" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"1D68" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"1D69" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"1D6A" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"1D6B" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"1D6C" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"1D6D" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"1D6E" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"1D6F" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"1D70" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"1D71" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"1D72" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"1D73" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"1D74" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"1D75" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"1D76" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"1D77" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"1D78" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"1D79" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"1D7A" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"1D7B" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"1D7C" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"1D7D" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"1D7E" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"1D7F" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"1D80" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"1D81" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"1D82" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"1D83" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"1D84" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"1D85" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"1D86" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"1D87" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"1D88" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"1D89" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"1D8A" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"1D8B" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"1D8C" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"1D8D" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"1D8E" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"1D8F" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"1D90" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"1D91" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"1D92" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"1D93" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"1D94" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"1D95" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"1D96" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"1D97" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"1D98" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"1D99" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"1D9A" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"1D9B" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"1D9C" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"1D9D" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"1D9E" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"1D9F" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"1DA0" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"1DA1" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"1DA2" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"1DA3" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"1DA4" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"1DA5" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"1DA6" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"1DA7" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"1DA8" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"1DA9" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"1DAA" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"1DAB" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"1DAC" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"1DAD" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"1DAE" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"1DAF" => MILLIEMES <= x"7"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"1DB0" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"1DB1" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"1DB2" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"1DB3" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"1DB4" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"1DB5" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"1DB6" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"1DB7" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"1DB8" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"1DB9" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"1DBA" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"1DBB" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"1DBC" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"1DBD" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"1DBE" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"1DBF" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"1DC0" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"1DC1" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"1DC2" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"1DC3" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"1DC4" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"1DC5" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"1DC6" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"1DC7" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"1DC8" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"1DC9" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"1DCA" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"1DCB" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"1DCC" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"1DCD" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"1DCE" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"1DCF" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"1DD0" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"1DD1" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"1DD2" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"1DD3" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"1DD4" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"1DD5" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"1DD6" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"1DD7" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"1DD8" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"1DD9" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"1DDA" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"1DDB" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"1DDC" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"1DDD" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"1DDE" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"1DDF" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"1DE0" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"1DE1" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"1DE2" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"1DE3" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"1DE4" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"1DE5" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"1DE6" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"1DE7" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"1DE8" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"1DE9" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"1DEA" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"1DEB" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"1DEC" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"1DED" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"1DEE" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"1DEF" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"1DF0" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"1DF1" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"1DF2" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"1DF3" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"1DF4" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"1DF5" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"1DF6" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"1DF7" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"1DF8" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"1DF9" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"1DFA" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"1DFB" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"1DFC" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"1DFD" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"1DFE" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"1DFF" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"1E00" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"1E01" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"1E02" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"1E03" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"1E04" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"1E05" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"1E06" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"1E07" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"1E08" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"1E09" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"1E0A" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"1E0B" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"1E0C" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"1E0D" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"1E0E" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"1E0F" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"1E10" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"1E11" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"1E12" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"1E13" => MILLIEMES <= x"7"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"1E14" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"1E15" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"1E16" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"1E17" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"1E18" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"1E19" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"1E1A" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"1E1B" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"1E1C" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"1E1D" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"1E1E" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"1E1F" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"1E20" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"1E21" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"1E22" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"1E23" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"1E24" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"1E25" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"1E26" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"1E27" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"1E28" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"1E29" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"1E2A" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"1E2B" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"1E2C" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"1E2D" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"1E2E" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"1E2F" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"1E30" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"1E31" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"1E32" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"1E33" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"1E34" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"1E35" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"1E36" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"1E37" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"1E38" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"1E39" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"1E3A" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"1E3B" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"1E3C" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"1E3D" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"1E3E" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"1E3F" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"1E40" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"1E41" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"1E42" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"1E43" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"1E44" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"1E45" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"1E46" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"1E47" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"1E48" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"1E49" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"1E4A" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"1E4B" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"1E4C" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"1E4D" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"1E4E" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"1E4F" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"1E50" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"1E51" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"1E52" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"1E53" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"1E54" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"1E55" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"1E56" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"1E57" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"1E58" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"1E59" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"1E5A" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"1E5B" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"1E5C" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"1E5D" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"1E5E" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"1E5F" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"1E60" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"1E61" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"1E62" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"1E63" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"1E64" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"1E65" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"1E66" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"1E67" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"1E68" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"1E69" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"1E6A" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"1E6B" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"1E6C" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"1E6D" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"1E6E" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"1E6F" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"1E70" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"1E71" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"1E72" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"1E73" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"1E74" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"1E75" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"1E76" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"1E77" => MILLIEMES <= x"7"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"1E78" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"1E79" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"1E7A" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"1E7B" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"1E7C" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"1E7D" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"1E7E" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"1E7F" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"1E80" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"1E81" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"1E82" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"1E83" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"1E84" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"1E85" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"1E86" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"1E87" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"1E88" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"1E89" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"1E8A" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"1E8B" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"1E8C" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"1E8D" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"1E8E" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"1E8F" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"1E90" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"1E91" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"1E92" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"1E93" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"1E94" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"1E95" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"1E96" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"1E97" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"1E98" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"1E99" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"1E9A" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"1E9B" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"1E9C" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"1E9D" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"1E9E" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"1E9F" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"1EA0" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"1EA1" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"1EA2" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"1EA3" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"1EA4" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"1EA5" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"1EA6" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"1EA7" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"1EA8" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"1EA9" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"1EAA" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"1EAB" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"1EAC" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"1EAD" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"1EAE" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"1EAF" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"1EB0" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"1EB1" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"1EB2" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"1EB3" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"1EB4" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"1EB5" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"1EB6" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"1EB7" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"1EB8" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"1EB9" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"1EBA" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"1EBB" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"1EBC" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"1EBD" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"1EBE" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"1EBF" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"1EC0" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"1EC1" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"1EC2" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"1EC3" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"1EC4" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"1EC5" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"1EC6" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"1EC7" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"1EC8" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"1EC9" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"1ECA" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"1ECB" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"1ECC" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"1ECD" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"1ECE" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"1ECF" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"1ED0" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"1ED1" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"1ED2" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"1ED3" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"1ED4" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"1ED5" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"1ED6" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"1ED7" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"1ED8" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"1ED9" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"1EDA" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"1EDB" => MILLIEMES <= x"7"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"1EDC" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"1EDD" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"1EDE" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"1EDF" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"1EE0" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"1EE1" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"1EE2" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"1EE3" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"1EE4" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"1EE5" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"1EE6" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"1EE7" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"1EE8" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"1EE9" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"1EEA" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"1EEB" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"1EEC" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"1EED" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"1EEE" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"1EEF" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"1EF0" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"1EF1" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"1EF2" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"1EF3" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"1EF4" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"1EF5" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"1EF6" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"1EF7" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"1EF8" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"1EF9" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"1EFA" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"1EFB" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"1EFC" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"1EFD" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"1EFE" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"1EFF" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"1F00" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"1F01" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"1F02" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"1F03" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"1F04" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"1F05" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"1F06" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"1F07" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"1F08" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"1F09" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"1F0A" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"1F0B" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"1F0C" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"1F0D" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"1F0E" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"1F0F" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"1F10" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"1F11" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"1F12" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"1F13" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"1F14" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"1F15" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"1F16" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"1F17" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"1F18" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"1F19" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"1F1A" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"1F1B" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"1F1C" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"1F1D" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"1F1E" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"1F1F" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"1F20" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"1F21" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"1F22" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"1F23" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"1F24" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"1F25" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"1F26" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"1F27" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"1F28" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"1F29" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"1F2A" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"1F2B" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"1F2C" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"1F2D" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"1F2E" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"1F2F" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"1F30" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"1F31" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"1F32" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"1F33" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"1F34" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"1F35" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"1F36" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"1F37" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"1F38" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"1F39" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"1F3A" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"1F3B" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"1F3C" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"1F3D" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"1F3E" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"1F3F" => MILLIEMES <= x"7"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"1F40" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"1F41" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"1F42" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"1F43" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"1F44" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"1F45" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"1F46" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"1F47" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"1F48" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"1F49" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"1F4A" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"1F4B" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"1F4C" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"1F4D" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"1F4E" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"1F4F" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"1F50" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"1F51" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"1F52" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"1F53" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"1F54" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"1F55" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"1F56" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"1F57" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"1F58" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"1F59" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"1F5A" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"1F5B" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"1F5C" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"1F5D" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"1F5E" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"1F5F" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"1F60" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"1F61" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"1F62" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"1F63" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"1F64" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"1F65" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"1F66" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"1F67" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"1F68" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"1F69" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"1F6A" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"1F6B" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"1F6C" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"1F6D" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"1F6E" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"1F6F" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"1F70" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"1F71" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"1F72" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"1F73" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"1F74" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"1F75" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"1F76" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"1F77" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"1F78" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"1F79" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"1F7A" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"1F7B" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"1F7C" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"1F7D" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"1F7E" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"1F7F" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"1F80" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"1F81" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"1F82" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"1F83" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"1F84" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"1F85" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"1F86" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"1F87" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"1F88" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"1F89" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"1F8A" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"1F8B" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"1F8C" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"1F8D" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"1F8E" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"1F8F" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"1F90" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"1F91" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"1F92" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"1F93" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"1F94" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"1F95" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"1F96" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"1F97" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"1F98" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"1F99" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"1F9A" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"1F9B" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"1F9C" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"1F9D" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"1F9E" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"1F9F" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"1FA0" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"1FA1" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"1FA2" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"1FA3" => MILLIEMES <= x"8"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"1FA4" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"1FA5" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"1FA6" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"1FA7" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"1FA8" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"1FA9" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"1FAA" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"1FAB" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"1FAC" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"1FAD" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"1FAE" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"1FAF" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"1FB0" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"1FB1" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"1FB2" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"1FB3" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"1FB4" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"1FB5" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"1FB6" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"1FB7" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"1FB8" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"1FB9" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"1FBA" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"1FBB" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"1FBC" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"1FBD" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"1FBE" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"1FBF" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"1FC0" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"1FC1" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"1FC2" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"1FC3" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"1FC4" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"1FC5" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"1FC6" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"1FC7" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"1FC8" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"1FC9" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"1FCA" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"1FCB" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"1FCC" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"1FCD" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"1FCE" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"1FCF" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"1FD0" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"1FD1" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"1FD2" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"1FD3" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"1FD4" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"1FD5" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"1FD6" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"1FD7" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"1FD8" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"1FD9" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"1FDA" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"1FDB" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"1FDC" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"1FDD" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"1FDE" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"1FDF" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"1FE0" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"1FE1" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"1FE2" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"1FE3" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"1FE4" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"1FE5" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"1FE6" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"1FE7" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"1FE8" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"1FE9" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"1FEA" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"1FEB" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"1FEC" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"1FED" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"1FEE" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"1FEF" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"1FF0" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"1FF1" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"1FF2" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"1FF3" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"1FF4" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"1FF5" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"1FF6" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"1FF7" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"1FF8" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"1FF9" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"1FFA" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"1FFB" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"1FFC" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"1FFD" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"1FFE" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"1FFF" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"2000" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"2001" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"2002" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"2003" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"2004" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"2005" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"2006" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"2007" => MILLIEMES <= x"8"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"2008" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"2009" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"200A" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"200B" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"200C" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"200D" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"200E" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"200F" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"2010" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"2011" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"2012" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"2013" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"2014" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"2015" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"2016" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"2017" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"2018" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"2019" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"201A" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"201B" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"201C" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"201D" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"201E" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"201F" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"2020" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"2021" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"2022" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"2023" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"2024" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"2025" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"2026" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"2027" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"2028" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"2029" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"202A" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"202B" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"202C" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"202D" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"202E" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"202F" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"2030" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"2031" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"2032" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"2033" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"2034" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"2035" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"2036" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"2037" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"2038" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"2039" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"203A" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"203B" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"203C" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"203D" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"203E" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"203F" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"2040" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"2041" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"2042" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"2043" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"2044" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"2045" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"2046" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"2047" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"2048" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"2049" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"204A" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"204B" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"204C" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"204D" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"204E" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"204F" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"2050" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"2051" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"2052" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"2053" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"2054" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"2055" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"2056" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"2057" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"2058" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"2059" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"205A" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"205B" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"205C" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"205D" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"205E" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"205F" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"2060" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"2061" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"2062" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"2063" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"2064" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"2065" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"2066" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"2067" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"2068" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"2069" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"206A" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"206B" => MILLIEMES <= x"8"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"206C" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"206D" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"206E" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"206F" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"2070" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"2071" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"2072" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"2073" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"2074" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"2075" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"2076" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"2077" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"2078" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"2079" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"207A" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"207B" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"207C" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"207D" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"207E" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"207F" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"2080" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"2081" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"2082" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"2083" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"2084" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"2085" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"2086" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"2087" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"2088" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"2089" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"208A" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"208B" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"208C" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"208D" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"208E" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"208F" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"2090" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"2091" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"2092" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"2093" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"2094" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"2095" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"2096" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"2097" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"2098" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"2099" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"209A" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"209B" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"209C" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"209D" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"209E" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"209F" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"20A0" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"20A1" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"20A2" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"20A3" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"20A4" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"20A5" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"20A6" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"20A7" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"20A8" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"20A9" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"20AA" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"20AB" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"20AC" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"20AD" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"20AE" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"20AF" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"20B0" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"20B1" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"20B2" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"20B3" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"20B4" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"20B5" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"20B6" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"20B7" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"20B8" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"20B9" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"20BA" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"20BB" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"20BC" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"20BD" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"20BE" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"20BF" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"20C0" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"20C1" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"20C2" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"20C3" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"20C4" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"20C5" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"20C6" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"20C7" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"20C8" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"20C9" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"20CA" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"20CB" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"20CC" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"20CD" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"20CE" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"20CF" => MILLIEMES <= x"8"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"20D0" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"20D1" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"20D2" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"20D3" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"20D4" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"20D5" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"20D6" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"20D7" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"20D8" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"20D9" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"20DA" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"20DB" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"20DC" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"20DD" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"20DE" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"20DF" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"20E0" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"20E1" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"20E2" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"20E3" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"20E4" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"20E5" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"20E6" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"20E7" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"20E8" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"20E9" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"20EA" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"20EB" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"20EC" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"20ED" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"20EE" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"20EF" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"20F0" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"20F1" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"20F2" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"20F3" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"20F4" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"20F5" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"20F6" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"20F7" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"20F8" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"20F9" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"20FA" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"20FB" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"20FC" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"20FD" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"20FE" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"20FF" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"2100" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"2101" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"2102" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"2103" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"2104" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"2105" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"2106" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"2107" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"2108" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"2109" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"210A" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"210B" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"210C" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"210D" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"210E" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"210F" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"2110" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"2111" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"2112" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"2113" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"2114" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"2115" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"2116" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"2117" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"2118" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"2119" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"211A" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"211B" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"211C" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"211D" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"211E" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"211F" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"2120" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"2121" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"2122" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"2123" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"2124" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"2125" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"2126" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"2127" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"2128" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"2129" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"212A" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"212B" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"212C" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"212D" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"212E" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"212F" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"2130" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"2131" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"2132" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"2133" => MILLIEMES <= x"8"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"2134" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"2135" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"2136" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"2137" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"2138" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"2139" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"213A" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"213B" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"213C" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"213D" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"213E" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"213F" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"2140" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"2141" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"2142" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"2143" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"2144" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"2145" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"2146" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"2147" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"2148" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"2149" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"214A" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"214B" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"214C" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"214D" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"214E" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"214F" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"2150" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"2151" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"2152" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"2153" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"2154" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"2155" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"2156" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"2157" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"2158" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"2159" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"215A" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"215B" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"215C" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"215D" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"215E" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"215F" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"2160" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"2161" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"2162" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"2163" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"2164" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"2165" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"2166" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"2167" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"2168" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"2169" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"216A" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"216B" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"216C" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"216D" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"216E" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"216F" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"2170" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"2171" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"2172" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"2173" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"2174" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"2175" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"2176" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"2177" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"2178" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"2179" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"217A" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"217B" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"217C" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"217D" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"217E" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"217F" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"2180" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"2181" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"2182" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"2183" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"2184" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"2185" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"2186" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"2187" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"2188" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"2189" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"218A" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"218B" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"218C" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"218D" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"218E" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"218F" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"2190" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"2191" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"2192" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"2193" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"2194" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"2195" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"2196" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"2197" => MILLIEMES <= x"8"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"2198" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"2199" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"219A" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"219B" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"219C" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"219D" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"219E" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"219F" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"21A0" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"21A1" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"21A2" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"21A3" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"21A4" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"21A5" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"21A6" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"21A7" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"21A8" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"21A9" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"21AA" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"21AB" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"21AC" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"21AD" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"21AE" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"21AF" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"21B0" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"21B1" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"21B2" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"21B3" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"21B4" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"21B5" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"21B6" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"21B7" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"21B8" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"21B9" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"21BA" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"21BB" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"21BC" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"21BD" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"21BE" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"21BF" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"21C0" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"21C1" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"21C2" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"21C3" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"21C4" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"21C5" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"21C6" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"21C7" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"21C8" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"21C9" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"21CA" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"21CB" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"21CC" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"21CD" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"21CE" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"21CF" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"21D0" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"21D1" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"21D2" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"21D3" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"21D4" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"21D5" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"21D6" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"21D7" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"21D8" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"21D9" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"21DA" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"21DB" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"21DC" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"21DD" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"21DE" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"21DF" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"21E0" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"21E1" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"21E2" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"21E3" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"21E4" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"21E5" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"21E6" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"21E7" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"21E8" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"21E9" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"21EA" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"21EB" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"21EC" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"21ED" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"21EE" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"21EF" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"21F0" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"21F1" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"21F2" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"21F3" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"21F4" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"21F5" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"21F6" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"21F7" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"21F8" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"21F9" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"21FA" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"21FB" => MILLIEMES <= x"8"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"21FC" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"21FD" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"21FE" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"21FF" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"2200" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"2201" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"2202" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"2203" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"2204" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"2205" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"2206" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"2207" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"2208" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"2209" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"220A" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"220B" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"220C" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"220D" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"220E" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"220F" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"2210" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"2211" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"2212" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"2213" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"2214" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"2215" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"2216" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"2217" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"2218" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"2219" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"221A" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"221B" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"221C" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"221D" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"221E" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"221F" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"2220" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"2221" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"2222" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"2223" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"2224" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"2225" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"2226" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"2227" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"2228" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"2229" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"222A" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"222B" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"222C" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"222D" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"222E" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"222F" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"2230" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"2231" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"2232" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"2233" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"2234" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"2235" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"2236" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"2237" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"2238" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"2239" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"223A" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"223B" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"223C" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"223D" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"223E" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"223F" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"2240" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"2241" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"2242" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"2243" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"2244" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"2245" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"2246" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"2247" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"2248" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"2249" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"224A" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"224B" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"224C" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"224D" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"224E" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"224F" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"2250" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"2251" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"2252" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"2253" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"2254" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"2255" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"2256" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"2257" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"2258" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"2259" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"225A" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"225B" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"225C" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"225D" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"225E" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"225F" => MILLIEMES <= x"8"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"2260" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"2261" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"2262" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"2263" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"2264" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"2265" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"2266" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"2267" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"2268" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"2269" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"226A" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"226B" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"226C" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"226D" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"226E" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"226F" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"2270" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"2271" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"2272" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"2273" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"2274" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"2275" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"2276" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"2277" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"2278" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"2279" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"227A" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"227B" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"227C" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"227D" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"227E" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"227F" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"2280" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"2281" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"2282" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"2283" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"2284" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"2285" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"2286" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"2287" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"2288" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"2289" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"228A" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"228B" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"228C" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"228D" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"228E" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"228F" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"2290" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"2291" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"2292" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"2293" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"2294" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"2295" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"2296" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"2297" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"2298" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"2299" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"229A" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"229B" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"229C" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"229D" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"229E" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"229F" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"22A0" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"22A1" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"22A2" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"22A3" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"22A4" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"22A5" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"22A6" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"22A7" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"22A8" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"22A9" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"22AA" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"22AB" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"22AC" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"22AD" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"22AE" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"22AF" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"22B0" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"22B1" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"22B2" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"22B3" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"22B4" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"22B5" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"22B6" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"22B7" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"22B8" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"22B9" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"22BA" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"22BB" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"22BC" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"22BD" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"22BE" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"22BF" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"22C0" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"22C1" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"22C2" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"22C3" => MILLIEMES <= x"8"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"22C4" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"22C5" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"22C6" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"22C7" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"22C8" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"22C9" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"22CA" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"22CB" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"22CC" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"22CD" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"22CE" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"22CF" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"22D0" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"22D1" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"22D2" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"22D3" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"22D4" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"22D5" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"22D6" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"22D7" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"22D8" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"22D9" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"22DA" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"22DB" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"22DC" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"22DD" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"22DE" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"22DF" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"22E0" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"22E1" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"22E2" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"22E3" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"22E4" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"22E5" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"22E6" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"22E7" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"22E8" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"22E9" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"22EA" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"22EB" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"22EC" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"22ED" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"22EE" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"22EF" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"22F0" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"22F1" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"22F2" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"22F3" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"22F4" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"22F5" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"22F6" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"22F7" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"22F8" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"22F9" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"22FA" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"22FB" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"22FC" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"22FD" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"22FE" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"22FF" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"2300" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"2301" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"2302" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"2303" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"2304" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"2305" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"2306" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"2307" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"2308" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"2309" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"230A" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"230B" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"230C" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"230D" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"230E" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"230F" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"2310" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"2311" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"2312" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"2313" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"2314" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"2315" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"2316" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"2317" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"2318" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"2319" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"231A" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"231B" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"231C" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"231D" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"231E" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"231F" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"2320" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"2321" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"2322" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"2323" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"2324" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"2325" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"2326" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"2327" => MILLIEMES <= x"8"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"2328" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"2329" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"232A" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"232B" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"232C" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"232D" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"232E" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"232F" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"2330" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"2331" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"2332" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"2333" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"2334" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"2335" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"2336" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"2337" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"2338" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"2339" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"233A" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"233B" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"233C" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"233D" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"233E" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"233F" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"2340" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"2341" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"2342" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"2343" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"2344" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"2345" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"2346" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"2347" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"2348" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"2349" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"234A" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"234B" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"234C" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"234D" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"234E" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"234F" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"2350" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"2351" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"2352" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"2353" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"2354" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"2355" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"2356" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"2357" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"2358" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"2359" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"235A" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"235B" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"235C" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"235D" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"235E" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"235F" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"2360" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"2361" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"2362" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"2363" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"2364" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"2365" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"2366" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"2367" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"2368" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"2369" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"236A" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"236B" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"236C" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"236D" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"236E" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"236F" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"2370" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"2371" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"2372" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"2373" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"2374" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"2375" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"2376" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"2377" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"2378" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"2379" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"237A" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"237B" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"237C" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"237D" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"237E" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"237F" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"2380" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"2381" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"2382" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"2383" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"2384" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"2385" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"2386" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"2387" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"2388" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"2389" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"238A" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"238B" => MILLIEMES <= x"9"; CENTAINES <= x"0"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"238C" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"238D" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"238E" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"238F" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"2390" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"2391" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"2392" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"2393" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"2394" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"2395" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"2396" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"2397" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"2398" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"2399" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"239A" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"239B" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"239C" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"239D" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"239E" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"239F" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"23A0" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"23A1" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"23A2" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"23A3" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"23A4" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"23A5" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"23A6" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"23A7" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"23A8" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"23A9" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"23AA" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"23AB" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"23AC" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"23AD" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"23AE" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"23AF" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"23B0" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"23B1" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"23B2" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"23B3" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"23B4" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"23B5" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"23B6" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"23B7" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"23B8" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"23B9" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"23BA" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"23BB" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"23BC" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"23BD" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"23BE" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"23BF" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"23C0" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"23C1" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"23C2" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"23C3" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"23C4" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"23C5" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"23C6" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"23C7" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"23C8" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"23C9" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"23CA" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"23CB" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"23CC" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"23CD" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"23CE" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"23CF" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"23D0" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"23D1" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"23D2" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"23D3" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"23D4" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"23D5" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"23D6" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"23D7" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"23D8" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"23D9" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"23DA" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"23DB" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"23DC" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"23DD" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"23DE" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"23DF" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"23E0" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"23E1" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"23E2" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"23E3" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"23E4" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"23E5" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"23E6" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"23E7" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"23E8" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"23E9" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"23EA" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"23EB" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"23EC" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"23ED" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"23EE" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"23EF" => MILLIEMES <= x"9"; CENTAINES <= x"1"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"23F0" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"23F1" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"23F2" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"23F3" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"23F4" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"23F5" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"23F6" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"23F7" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"23F8" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"23F9" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"23FA" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"23FB" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"23FC" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"23FD" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"23FE" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"23FF" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"2400" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"2401" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"2402" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"2403" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"2404" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"2405" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"2406" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"2407" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"2408" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"2409" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"240A" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"240B" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"240C" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"240D" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"240E" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"240F" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"2410" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"2411" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"2412" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"2413" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"2414" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"2415" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"2416" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"2417" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"2418" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"2419" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"241A" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"241B" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"241C" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"241D" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"241E" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"241F" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"2420" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"2421" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"2422" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"2423" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"2424" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"2425" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"2426" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"2427" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"2428" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"2429" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"242A" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"242B" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"242C" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"242D" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"242E" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"242F" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"2430" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"2431" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"2432" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"2433" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"2434" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"2435" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"2436" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"2437" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"2438" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"2439" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"243A" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"243B" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"243C" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"243D" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"243E" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"243F" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"2440" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"2441" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"2442" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"2443" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"2444" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"2445" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"2446" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"2447" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"2448" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"2449" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"244A" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"244B" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"244C" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"244D" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"244E" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"244F" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"2450" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"2451" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"2452" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"2453" => MILLIEMES <= x"9"; CENTAINES <= x"2"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"2454" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"2455" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"2456" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"2457" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"2458" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"2459" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"245A" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"245B" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"245C" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"245D" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"245E" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"245F" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"2460" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"2461" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"2462" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"2463" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"2464" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"2465" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"2466" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"2467" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"2468" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"2469" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"246A" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"246B" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"246C" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"246D" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"246E" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"246F" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"2470" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"2471" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"2472" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"2473" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"2474" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"2475" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"2476" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"2477" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"2478" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"2479" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"247A" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"247B" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"247C" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"247D" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"247E" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"247F" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"2480" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"2481" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"2482" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"2483" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"2484" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"2485" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"2486" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"2487" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"2488" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"2489" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"248A" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"248B" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"248C" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"248D" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"248E" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"248F" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"2490" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"2491" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"2492" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"2493" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"2494" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"2495" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"2496" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"2497" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"2498" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"2499" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"249A" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"249B" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"249C" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"249D" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"249E" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"249F" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"24A0" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"24A1" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"24A2" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"24A3" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"24A4" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"24A5" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"24A6" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"24A7" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"24A8" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"24A9" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"24AA" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"24AB" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"24AC" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"24AD" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"24AE" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"24AF" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"24B0" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"24B1" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"24B2" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"24B3" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"24B4" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"24B5" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"24B6" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"24B7" => MILLIEMES <= x"9"; CENTAINES <= x"3"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"24B8" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"24B9" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"24BA" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"24BB" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"24BC" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"24BD" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"24BE" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"24BF" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"24C0" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"24C1" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"24C2" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"24C3" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"24C4" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"24C5" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"24C6" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"24C7" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"24C8" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"24C9" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"24CA" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"24CB" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"24CC" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"24CD" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"24CE" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"24CF" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"24D0" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"24D1" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"24D2" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"24D3" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"24D4" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"24D5" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"24D6" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"24D7" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"24D8" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"24D9" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"24DA" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"24DB" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"24DC" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"24DD" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"24DE" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"24DF" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"24E0" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"24E1" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"24E2" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"24E3" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"24E4" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"24E5" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"24E6" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"24E7" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"24E8" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"24E9" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"24EA" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"24EB" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"24EC" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"24ED" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"24EE" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"24EF" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"24F0" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"24F1" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"24F2" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"24F3" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"24F4" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"24F5" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"24F6" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"24F7" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"24F8" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"24F9" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"24FA" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"24FB" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"24FC" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"24FD" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"24FE" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"24FF" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"2500" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"2501" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"2502" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"2503" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"2504" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"2505" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"2506" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"2507" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"2508" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"2509" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"250A" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"250B" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"250C" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"250D" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"250E" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"250F" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"2510" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"2511" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"2512" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"2513" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"2514" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"2515" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"2516" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"2517" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"2518" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"2519" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"251A" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"251B" => MILLIEMES <= x"9"; CENTAINES <= x"4"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"251C" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"251D" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"251E" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"251F" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"2520" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"2521" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"2522" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"2523" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"2524" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"2525" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"2526" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"2527" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"2528" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"2529" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"252A" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"252B" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"252C" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"252D" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"252E" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"252F" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"2530" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"2531" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"2532" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"2533" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"2534" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"2535" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"2536" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"2537" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"2538" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"2539" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"253A" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"253B" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"253C" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"253D" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"253E" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"253F" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"2540" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"2541" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"2542" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"2543" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"2544" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"2545" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"2546" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"2547" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"2548" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"2549" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"254A" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"254B" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"254C" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"254D" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"254E" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"254F" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"2550" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"2551" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"2552" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"2553" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"2554" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"2555" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"2556" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"2557" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"2558" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"2559" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"255A" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"255B" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"255C" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"255D" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"255E" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"255F" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"2560" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"2561" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"2562" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"2563" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"2564" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"2565" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"2566" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"2567" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"2568" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"2569" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"256A" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"256B" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"256C" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"256D" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"256E" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"256F" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"2570" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"2571" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"2572" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"2573" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"2574" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"2575" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"2576" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"2577" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"2578" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"2579" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"257A" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"257B" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"257C" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"257D" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"257E" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"257F" => MILLIEMES <= x"9"; CENTAINES <= x"5"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"2580" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"2581" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"2582" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"2583" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"2584" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"2585" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"2586" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"2587" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"2588" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"2589" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"258A" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"258B" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"258C" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"258D" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"258E" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"258F" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"2590" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"2591" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"2592" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"2593" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"2594" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"2595" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"2596" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"2597" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"2598" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"2599" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"259A" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"259B" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"259C" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"259D" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"259E" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"259F" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"25A0" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"25A1" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"25A2" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"25A3" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"25A4" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"25A5" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"25A6" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"25A7" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"25A8" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"25A9" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"25AA" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"25AB" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"25AC" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"25AD" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"25AE" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"25AF" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"25B0" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"25B1" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"25B2" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"25B3" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"25B4" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"25B5" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"25B6" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"25B7" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"25B8" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"25B9" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"25BA" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"25BB" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"25BC" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"25BD" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"25BE" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"25BF" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"25C0" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"25C1" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"25C2" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"25C3" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"25C4" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"25C5" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"25C6" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"25C7" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"25C8" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"25C9" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"25CA" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"25CB" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"25CC" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"25CD" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"25CE" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"25CF" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"25D0" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"25D1" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"25D2" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"25D3" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"25D4" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"25D5" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"25D6" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"25D7" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"25D8" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"25D9" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"25DA" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"25DB" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"25DC" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"25DD" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"25DE" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"25DF" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"25E0" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"25E1" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"25E2" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"25E3" => MILLIEMES <= x"9"; CENTAINES <= x"6"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"25E4" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"25E5" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"25E6" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"25E7" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"25E8" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"25E9" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"25EA" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"25EB" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"25EC" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"25ED" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"25EE" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"25EF" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"25F0" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"25F1" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"25F2" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"25F3" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"25F4" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"25F5" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"25F6" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"25F7" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"25F8" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"25F9" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"25FA" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"25FB" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"25FC" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"25FD" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"25FE" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"25FF" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"2600" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"2601" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"2602" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"2603" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"2604" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"2605" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"2606" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"2607" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"2608" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"2609" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"260A" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"260B" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"260C" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"260D" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"260E" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"260F" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"2610" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"2611" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"2612" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"2613" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"2614" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"2615" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"2616" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"2617" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"2618" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"2619" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"261A" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"261B" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"261C" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"261D" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"261E" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"261F" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"2620" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"2621" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"2622" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"2623" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"2624" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"2625" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"2626" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"2627" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"2628" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"2629" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"262A" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"262B" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"262C" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"262D" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"262E" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"262F" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"2630" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"2631" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"2632" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"2633" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"2634" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"2635" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"2636" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"2637" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"2638" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"2639" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"263A" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"263B" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"263C" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"263D" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"263E" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"263F" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"2640" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"2641" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"2642" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"2643" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"2644" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"2645" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"2646" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"2647" => MILLIEMES <= x"9"; CENTAINES <= x"7"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"2648" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"2649" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"264A" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"264B" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"264C" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"264D" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"264E" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"264F" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"2650" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"2651" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"2652" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"2653" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"2654" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"2655" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"2656" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"2657" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"2658" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"2659" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"265A" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"265B" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"265C" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"265D" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"265E" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"265F" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"2660" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"2661" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"2662" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"2663" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"2664" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"2665" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"2666" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"2667" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"2668" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"2669" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"266A" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"266B" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"266C" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"266D" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"266E" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"266F" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"2670" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"2671" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"2672" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"2673" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"2674" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"2675" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"2676" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"2677" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"2678" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"2679" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"267A" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"267B" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"267C" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"267D" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"267E" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"267F" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"2680" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"2681" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"2682" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"2683" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"2684" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"2685" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"2686" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"2687" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"2688" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"2689" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"268A" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"268B" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"268C" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"268D" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"268E" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"268F" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"2690" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"2691" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"2692" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"2693" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"2694" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"2695" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"2696" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"2697" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"2698" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"2699" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"269A" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"269B" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"269C" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"269D" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"269E" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"269F" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"26A0" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"26A1" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"26A2" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"26A3" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"26A4" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"26A5" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"26A6" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"26A7" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"26A8" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"26A9" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"26AA" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"26AB" => MILLIEMES <= x"9"; CENTAINES <= x"8"; DIZAINES <= x"9"; UNITES <= x"9";
--			when x"26AC" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"0";
--			when x"26AD" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"1";
--			when x"26AE" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"2";
--			when x"26AF" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"3";
--			when x"26B0" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"4";
--			when x"26B1" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"5";
--			when x"26B2" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"6";
--			when x"26B3" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"7";
--			when x"26B4" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"8";
--			when x"26B5" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"0"; UNITES <= x"9";
--			when x"26B6" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"0";
--			when x"26B7" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"1";
--			when x"26B8" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"2";
--			when x"26B9" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"3";
--			when x"26BA" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"4";
--			when x"26BB" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"5";
--			when x"26BC" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"6";
--			when x"26BD" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"7";
--			when x"26BE" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"8";
--			when x"26BF" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"1"; UNITES <= x"9";
--			when x"26C0" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"0";
--			when x"26C1" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"1";
--			when x"26C2" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"2";
--			when x"26C3" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"3";
--			when x"26C4" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"4";
--			when x"26C5" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"5";
--			when x"26C6" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"6";
--			when x"26C7" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"7";
--			when x"26C8" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"8";
--			when x"26C9" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"2"; UNITES <= x"9";
--			when x"26CA" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"0";
--			when x"26CB" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"1";
--			when x"26CC" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"2";
--			when x"26CD" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"3";
--			when x"26CE" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"4";
--			when x"26CF" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"5";
--			when x"26D0" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"6";
--			when x"26D1" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"7";
--			when x"26D2" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"8";
--			when x"26D3" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"3"; UNITES <= x"9";
--			when x"26D4" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"0";
--			when x"26D5" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"1";
--			when x"26D6" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"2";
--			when x"26D7" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"3";
--			when x"26D8" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"4";
--			when x"26D9" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"5";
--			when x"26DA" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"6";
--			when x"26DB" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"7";
--			when x"26DC" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"8";
--			when x"26DD" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"4"; UNITES <= x"9";
--			when x"26DE" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"0";
--			when x"26DF" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"1";
--			when x"26E0" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"2";
--			when x"26E1" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"3";
--			when x"26E2" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"4";
--			when x"26E3" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"5";
--			when x"26E4" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"6";
--			when x"26E5" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"7";
--			when x"26E6" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"8";
--			when x"26E7" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"5"; UNITES <= x"9";
--			when x"26E8" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"0";
--			when x"26E9" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"1";
--			when x"26EA" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"2";
--			when x"26EB" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"3";
--			when x"26EC" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"4";
--			when x"26ED" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"5";
--			when x"26EE" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"6";
--			when x"26EF" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"7";
--			when x"26F0" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"8";
--			when x"26F1" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"6"; UNITES <= x"9";
--			when x"26F2" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"0";
--			when x"26F3" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"1";
--			when x"26F4" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"2";
--			when x"26F5" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"3";
--			when x"26F6" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"4";
--			when x"26F7" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"5";
--			when x"26F8" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"6";
--			when x"26F9" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"7";
--			when x"26FA" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"8";
--			when x"26FB" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"7"; UNITES <= x"9";
--			when x"26FC" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"0";
--			when x"26FD" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"1";
--			when x"26FE" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"2";
--			when x"26FF" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"3";
--			when x"2700" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"4";
--			when x"2701" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"5";
--			when x"2702" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"6";
--			when x"2703" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"7";
--			when x"2704" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"8";
--			when x"2705" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"8"; UNITES <= x"9";
--			when x"2706" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"0";
--			when x"2707" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"1";
--			when x"2708" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"2";
--			when x"2709" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"3";
--			when x"270A" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"4";
--			when x"270B" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"5";
--			when x"270C" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"6";
--			when x"270D" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"7";
--			when x"270E" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"8";
--			when x"270F" => MILLIEMES <= x"9"; CENTAINES <= x"9"; DIZAINES <= x"9"; UNITES <= x"9";
